module top_eco(\a[0] , n_506,\a[5] ,\b[2] ,\b[4] ,\b[5] ,\op[1] , n_505, n_474, wc1, n_482, wc3, n_489, n_490, wc7, n_495, wc17, n_504, wc20, n_508, wc21, n_480, wc22, n_488, wc52, wc26, n_492, wc27, wc42, wc61, overflow,\y[6] ,\y[7] ,\y[0] ,\y[1] ,\y[2] ,\y[3] ,\y[4] ,\y[5] , n_803, n_804);
  input \a[0] , n_506,\a[5] ,\b[2] ;
  input \b[4] ,\b[5] ,\op[1] , n_505, n_474;
  input wc1, n_482, wc3, n_489, n_490;
  input wc7, n_495, wc17, n_504, wc20;
  input n_508, wc21, n_480, wc22, n_488;
  input wc52, wc26, n_492, wc27, wc42;
  input wc61;
  output overflow,\y[6] ,\y[7] ,\y[0] ;
  output \y[1] ,\y[2] ,\y[3] ,\y[4] ,\y[5] ;
  output n_803, n_804;
  wire patchNew_n_264, patchNew_n_475, patchNew_n_496, patchNew_n_451;
  wire patchNew_wc10, patchNew_n_502, patchNew_n_804, patchNew_wc12, patchNew_n_450;
  wire patchNew_n_806, patchNew_n_805, patchNew_wc13, patchNew_n_807, patchNew_n_503;
  wire patchNew_n_811, patchNew_wc17, patchNew_n_812, patchNew_n_69, patchNew_n_505;
  wire patchNew_n_455, patchNew_n_705, patchNew_n_819, patchNew_n_820, patchNew_n_413;
  wire patchNew_n_522, patchNew_n_687, patchNew_n_369, patchNew_n_657, patchNew_n_410;
  wire patchNew_n_521, patchNew_n_615, patchNew_n_360, patchNew_n_579, patchNew_wc63;
  wire patchNew_wc66, patchNew_wc65, patchNew_wc68, patchNew_wc67, patchNew_wc69;
  and eco1 (\y[0] , n_495, patchNew_wc66);
  and eco2 (\y[1] , n_508, patchNew_wc63);
  and eco3 (\y[2] , n_480, patchNew_wc68);
  and eco4 (\y[3] , n_492, patchNew_wc67);
  and eco5 (\y[4] , n_488, patchNew_wc65);
  and eco6 (\y[5] , patchNew_wc69, n_504);
  or eco7 (n_803, patchNew_wc10, n_495);
  or eco8 (n_804, patchNew_n_451, wc17);
  assign overflow = \y[7] ;
  assign \y[6]  = \y[7] ;
  not eco11 (\y[7] , patchNew_n_69);
  nand eco12 (patchNew_n_451, patchNew_n_804, patchNew_n_805);
  not eco13 (patchNew_wc10, patchNew_n_451);
  nand eco14 (patchNew_n_502, patchNew_n_806, patchNew_n_807);
  or eco15 (patchNew_n_804, patchNew_wc12, patchNew_n_450);
  not eco16 (patchNew_wc12, patchNew_n_502);
  nand eco17 (patchNew_n_450, patchNew_n_811, patchNew_n_812);
  or eco18 (patchNew_n_806, wc20, n_480);
  or eco19 (patchNew_n_805, patchNew_n_502, patchNew_wc13);
  not eco20 (patchNew_wc13, patchNew_n_450);
  or eco21 (patchNew_n_807, n_504, wc22);
  nand eco22 (patchNew_n_503, patchNew_n_819, patchNew_n_820);
  or eco23 (patchNew_n_811, patchNew_wc17, n_488);
  not eco24 (patchNew_wc17, patchNew_n_503);
  or eco25 (patchNew_n_812, patchNew_n_503, wc26);
  or eco26 (patchNew_n_69, patchNew_n_505, patchNew_n_264);
  or eco27 (patchNew_n_819, wc27, n_508);
  or eco28 (patchNew_n_820, n_492, wc21);
  not eco29 (patchNew_wc63, patchNew_n_69);
  not eco30 (patchNew_wc66, patchNew_n_69);
  not eco31 (patchNew_wc65, patchNew_n_69);
  not eco32 (patchNew_wc68, patchNew_n_69);
  not eco33 (patchNew_wc67, patchNew_n_69);
  not eco34 (patchNew_wc69, patchNew_n_69);
  nand eco35 (patchNew_n_505, patchNew_n_455, patchNew_n_705);
  or eco36 (patchNew_n_264, wc52,\op[1] );
  or eco37 (patchNew_n_455, wc7,\b[5] );
  nand eco38 (patchNew_n_705, patchNew_n_475, patchNew_n_413);
  or eco39 (patchNew_n_475, wc61,\a[5] );
  nand eco40 (patchNew_n_413, patchNew_n_522, patchNew_n_687);
  or eco41 (patchNew_n_522, wc3,\b[4] );
  nand eco42 (patchNew_n_687, n_482, patchNew_n_369);
  nand eco43 (patchNew_n_369, n_490, patchNew_n_657);
  nand eco44 (patchNew_n_657, n_489, patchNew_n_410);
  nand eco45 (patchNew_n_410, patchNew_n_521, patchNew_n_615);
  or eco46 (patchNew_n_521, wc1,\b[2] );
  nand eco47 (patchNew_n_615, n_474, patchNew_n_360);
  nand eco48 (patchNew_n_360, n_506, patchNew_n_579);
  nand eco49 (patchNew_n_579, n_505, patchNew_n_496);
  or eco50 (patchNew_n_496, wc42,\a[0] );
endmodule
