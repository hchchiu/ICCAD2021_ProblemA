module top_eco(g4671, g4672, g4669, g4705, g4706, g4707, g4708, g4674, g4676, g4677, g4680, g4681, g4682, g4683, g4684, g4685, g4687, g4688, g4689, g4691, g4692, g4693, g4694, g4695, g4696, g4697, g4698, g4699, g4700, g4701, g4703, g4704, g471, g4709, g4710, g4711, g4715, g4716, g4717, g4718, g4719, g4720, g4721, g4725, g4726, g4727, g4729, g4731, g4732, g4735, g4736, g4738, g4740, g4741, g4743, g4744, g4746, g4748, g4749, g4750, g4751, g4752, g4753, g4754, g4755, g4756, g4757, g4758, g4764, g4766, g4767, g4768, g4769, g4770, g4771, g4772, g4773, g4774, g4775, g4776, g4778, g4779, g4780, g4781, g4782, g4784, g4785, g4787, g4788, g4789, g4790, g4791, g4793, g4794, g4795, g4796, g4797, g4798, g4799, g4800, g4802, g4803, g4806, g4807, g4808, g4809, g4810, g4811, g4812, g4813, g4814, g4815, g1357, g1240, g923, g445, g448, g450, g454, g460, g461, g476, g478, g483, g487, g491, g492, g495, g497, g501, g505, g509, g510, g511_g4785, g518, g533, g535, g536, g538, g542, g550, g553, g555, g569, g575, g576, g580, g581, g582, g593, g600, g608, g609, g610, g618, g624, g625, g627, g630, g632, g633, g643, g648, g658, g665, g670, g685, g686, g687, g688, g703, g705, g706, g710, g720, g724, g730, g731, g739, g750, g753, g760, g771, g790, g801, g804, g813, g839, g864, g878, g904, g953, g987, g1015, g1024, g1035, g1049, g4702_g4785, g1062, g1068, g1122, g1123, g1156, g1171, g1308, g1332, g1340, g4849, g4851, g4852, g4853, g4854, g4855, g4856, g4857, g4861, g4862, g4863, g4864, g4865, g4866, g4867, g4868, g4869, g4870, g4871, g4873, g4874, g4879, g4880, g4881, g4882, g4883, g4884, g4886, g4888, g4889, g992, g1350, g1358, g991, g983, g1352, g989, g1343, g1325, g1339);
  input g4671, g4672, g4669, g4705;
  input g4706, g4707, g4708, g4674, g4676;
  input g4677, g4680, g4681, g4682, g4683;
  input g4684, g4685, g4687, g4688, g4689;
  input g4691, g4692, g4693, g4694, g4695;
  input g4696, g4697, g4698, g4699, g4700;
  input g4701, g4703, g4704, g471, g4709;
  input g4710, g4711, g4715, g4716, g4717;
  input g4718, g4719, g4720, g4721, g4725;
  input g4726, g4727, g4729, g4731, g4732;
  input g4735, g4736, g4738, g4740, g4741;
  input g4743, g4744, g4746, g4748, g4749;
  input g4750, g4751, g4752, g4753, g4754;
  input g4755, g4756, g4757, g4758, g4764;
  input g4766, g4767, g4768, g4769, g4770;
  input g4771, g4772, g4773, g4774, g4775;
  input g4776, g4778, g4779, g4780, g4781;
  input g4782, g4784, g4785, g4787, g4788;
  input g4789, g4790, g4791, g4793, g4794;
  input g4795, g4796, g4797, g4798, g4799;
  input g4800, g4802, g4803, g4806, g4807;
  input g4808, g4809, g4810, g4811, g4812;
  input g4813, g4814, g4815, g1357, g1240;
  input g923, g445, g448, g450, g454;
  input g460, g461, g476, g478, g483;
  input g487, g491, g492, g495, g497;
  input g501, g505, g509, g510, g511_g4785;
  input g518, g533, g535, g536, g538;
  input g542, g550, g553, g555, g569;
  input g575, g576, g580, g581, g582;
  input g593, g600, g608, g609, g610;
  input g618, g624, g625, g627, g630;
  input g632, g633, g643, g648, g658;
  input g665, g670, g685, g686, g687;
  input g688, g703, g705, g706, g710;
  input g720, g724, g730, g731, g739;
  input g750, g753, g760, g771, g790;
  input g801, g804, g813, g839, g864;
  input g878, g904, g953, g987, g1015;
  input g1024, g1035, g1049, g4702_g4785, g1062;
  input g1068, g1122, g1123, g1156, g1171;
  input g1308, g1332, g1340;
  output g4849, g4851, g4852, g4853;
  output g4854, g4855, g4856, g4857, g4861;
  output g4862, g4863, g4864, g4865, g4866;
  output g4867, g4868, g4869, g4870, g4871;
  output g4873, g4874, g4879, g4880, g4881;
  output g4882, g4883, g4884, g4886, g4888;
  output g4889, g992, g1350, g1358, g991;
  output g983, g1352, g989, g1343, g1325;
  output g1339;
  buf eco1 (g4849, patchNew_n1040);
  buf eco2 (g4851, patchNew_n593);
  buf eco3 (g4852, patchNew_n477);
  buf eco4 (g4853, patchNew_n1037);
  buf eco5 (g4854, patchNew_n747);
  buf eco6 (g4855, patchNew_n770);
  buf eco7 (g4856, patchNew_n1031);
  buf eco8 (g4857, patchNew_n373);
  buf eco9 (g4861, patchNew_n244);
  buf eco10 (g4862, patchNew_n378);
  buf eco11 (g4863, patchNew_n1034);
  buf eco12 (g4864, patchNew_n400);
  buf eco13 (g4865, patchNew_n348);
  buf eco14 (g4866, patchNew_n448);
  buf eco15 (g4867, patchNew_n494);
  buf eco16 (g4868, patchNew_n1029);
  buf eco17 (g4869, patchNew_n1029);
  buf eco18 (g4870, patchNew_n1033);
  buf eco19 (g4871, patchNew_n1033);
  buf eco20 (g4873, patchNew_n1026);
  buf eco21 (g4874, patchNew_n1026);
  buf eco22 (g4879, patchNew_n976);
  buf eco23 (g4880, patchNew_n977);
  buf eco24 (g4881, patchNew_n1017);
  buf eco25 (g4882, patchNew_n1001);
  buf eco26 (g4883, patchNew_n1000);
  buf eco27 (g4884, patchNew_n1000);
  buf eco28 (g4886, patchNew_n588);
  buf eco29 (g4888, patchNew_n837);
  buf eco30 (g4889, patchNew_n838);
  nand eco31 (g992, patchNew_n139_n140_n141, g4810);
  nand eco32 (g1350, patchNew_n1043, g4787);
  nand eco33 (g1358, patchNew_n1045, g4815);
  not eco34 (g991, patchNew_n1040);
  nand eco35 (g983, g4790, patchNew_n321);
  nand eco36 (g1352, patchNew_n116_n121_n28, patchNew_n593);
  nand eco37 (g989, patchNew_n121_n1038_n116, patchNew_n593);
  nand eco38 (g1343, patchNew_n1021, patchNew_n1022);
  nand eco39 (g1325, patchNew_1'b1_n1018, patchNew__xnor_GATE_0);
  not eco40 (g1339, patchNew_n835);
  and eco41 (patchNew_n1040, patchNew_new_n263_, patchNew_new_n266_);
  nor eco42 (patchNew_n593, patchNew_new_n268_, patchNew_new_n269_);
  nor eco43 (patchNew_n1031, patchNew_new_n313_, patchNew_new_n314_);
  and eco44 (patchNew_n373, patchNew__not_GATE_23, patchNew_new_n324_);
  or eco45 (patchNew_n244, patchNew_new_n328_, patchNew__not_GATE_27);
  or eco46 (patchNew_n378, patchNew_new_n323_, patchNew_new_n333_);
  not eco47 (patchNew_n1034, patchNew_n1031);
  not eco48 (patchNew_n400, );
  or eco49 (patchNew_n448, patchNew_new_n344_, patchNew__not_GATE_32);
  or eco50 (patchNew_n1029, patchNew_new_n365_, patchNew_new_n366_);
  or eco51 (patchNew_n1033, patchNew_new_n368_, patchNew_new_n369_);
  or eco52 (patchNew_n1026, patchNew_new_n372_, patchNew_new_n382_);
  and eco53 (patchNew_n976, patchNew__not_GATE_86, patchNew_new_n532_);
  not eco54 (patchNew_n977, patchNew_n976);
  nor eco55 (patchNew_n1017, patchNew_new_n548_, patchNew_new_n551_);
  and eco56 (patchNew_n1001, patchNew__not_GATE_110, patchNew_new_n583_);
  or eco57 (patchNew_n1000, patchNew_new_n585_, patchNew_new_n609_);
  or eco58 (patchNew_n588, patchNew_new_n638_, patchNew_new_n701_);
  and eco59 (patchNew_n837, patchNew__not_GATE_179, patchNew_new_n721_);
  not eco60 (patchNew_n838, patchNew_n837);
  and eco61 (patchNew_n321, patchNew__not_GATE_41, patchNew_new_n380_);
  and eco62 (patchNew_new_n320_, g670, patchNew__not_GATE_21);
  or eco63 (patchNew_n835, patchNew_new_n715_, patchNew__not_GATE_177);
  buf eco64 (patchNew_1'b1_n1018, g4812);
  or eco65 (patchNew_n1021, g4790, patchNew_new_n371_);
  or eco66 (patchNew_n1022, g864, patchNew_new_n364_);
  nand eco67 (patchNew_n116_n121_n28, g987, g4696);
  or eco68 (patchNew_n121_n1038_n116, patchNew__not_GATE_183, patchNew_new_n730_);
  not eco69 (patchNew_n1043, g1357);
  buf eco70 (patchNew_n1045, patchNew_n1043);
  or eco71 (patchNew_n139_n140_n141, patchNew__not_GATE_184, patchNew_new_n732_);
  not eco72 (patchNew_n1050, g706);
  xnor eco73 (patchNew__xnor_GATE_4, patchNew_new_n587_, patchNew_new_n593_);
  xnor eco74 (patchNew__xnor_GATE_5, patchNew_n348, patchNew_n494);
  xnor eco75 (patchNew__xnor_GATE_6, g4809, patchNew_new_n486_);
  xnor eco76 (patchNew__xnor_GATE_7, g4793, patchNew_new_n493_);
  xnor eco77 (patchNew__xnor_GATE_8, patchNew_n477, patchNew_n1037);
  xnor eco78 (patchNew__xnor_GATE_9, patchNew_new_n371_, patchNew_new_n535_);
  xnor eco79 (patchNew__xnor_GATE_10, patchNew_n770, patchNew_new_n659_);
  xnor eco80 (patchNew__xnor_GATE_11, patchNew_new_n705_, patchNew_new_n710_);
  not eco81 (patchNew__not_GATE_100, patchNew_new_n413_);
  not eco82 (patchNew__not_GATE_101, patchNew_n747);
  and eco83 (patchNew_new_n562_, g1122, g4752);
  and eco84 (patchNew_new_n563_, g4782, g501);
  and eco85 (patchNew_new_n564_, g4772, g706);
  and eco86 (patchNew_new_n565_, patchNew__not_GATE_102, g497);
  not eco87 (patchNew__not_GATE_102, g1156);
  nor eco88 (patchNew_new_n566_, patchNew_new_n563_, patchNew_new_n564_);
  and eco89 (patchNew_new_n567_, patchNew__not_GATE_103, patchNew_new_n566_);
  not eco90 (patchNew__not_GATE_103, patchNew_new_n565_);
  nor eco91 (patchNew_new_n568_, patchNew_new_n562_, patchNew_new_n567_);
  not eco92 (patchNew__not_GATE_104, patchNew_new_n391_);
  not eco93 (patchNew__not_GATE_105, patchNew_new_n401_);
  and eco94 (patchNew_new_n572_, patchNew_new_n568_, patchNew__xnor_GATE_2);
  nor eco95 (patchNew_new_n573_, patchNew_new_n568_, patchNew__xnor_GATE_2);
  not eco96 (patchNew__not_GATE_106, patchNew_new_n574_);
  not eco97 (patchNew__not_GATE_107, patchNew_new_n511_);
  and eco98 (patchNew_new_n578_, patchNew__xnor_GATE_1, patchNew__xnor_GATE_3);
  nor eco99 (patchNew_new_n579_, patchNew__xnor_GATE_1, patchNew__xnor_GATE_3);
  nor eco100 (patchNew_new_n580_, patchNew_new_n578_, patchNew_new_n579_);
  and eco101 (patchNew_new_n581_, patchNew__not_GATE_108, patchNew_new_n580_);
  not eco102 (patchNew__not_GATE_108, patchNew_new_n558_);
  and eco103 (patchNew_new_n582_, patchNew_new_n558_, patchNew__not_GATE_109);
  not eco104 (patchNew__not_GATE_109, patchNew_new_n580_);
  nor eco105 (patchNew_new_n583_, g4697, patchNew_new_n581_);
  not eco106 (patchNew__not_GATE_110, patchNew_new_n582_);
  nor eco107 (patchNew_new_n585_, g4791, patchNew_new_n547_);
  and eco108 (patchNew_new_n586_, patchNew__not_GATE_111, patchNew_new_n547_);
  not eco109 (patchNew__not_GATE_111, patchNew_new_n490_);
  and eco110 (patchNew_new_n588_, patchNew_n244, patchNew_new_n371_);
  and eco111 (patchNew_new_n589_, patchNew_n244, patchNew_new_n364_);
  nor eco112 (patchNew_new_n590_, patchNew_n244, patchNew_new_n364_);
  nor eco113 (patchNew_new_n591_, patchNew_new_n589_, patchNew_new_n590_);
  and eco114 (patchNew_new_n592_, patchNew__not_GATE_112, patchNew_new_n591_);
  not eco115 (patchNew__not_GATE_112, patchNew_new_n371_);
  not eco116 (patchNew__not_GATE_113, patchNew_new_n593_);
  not eco117 (patchNew__not_GATE_114, patchNew_new_n587_);
  and eco118 (patchNew_new_n597_, patchNew_n770, patchNew_n448);
  nor eco119 (patchNew_new_n598_, patchNew_n770, patchNew_n448);
  nor eco120 (patchNew_new_n599_, patchNew_new_n597_, patchNew_new_n598_);
  not eco121 (patchNew__not_GATE_115, patchNew_n348);
  not eco122 (patchNew__not_GATE_116, patchNew_n494);
  and eco123 (patchNew_new_n603_, patchNew_new_n599_, patchNew__xnor_GATE_5);
  nor eco124 (patchNew_new_n604_, patchNew_new_n599_, patchNew__xnor_GATE_5);
  nor eco125 (patchNew_new_n605_, patchNew_new_n603_, patchNew_new_n604_);
  and eco126 (patchNew_new_n606_, patchNew__not_GATE_117, patchNew_new_n605_);
  not eco127 (patchNew__not_GATE_117, patchNew__xnor_GATE_4);
  and eco128 (patchNew_new_n607_, patchNew__not_GATE_118, patchNew__xnor_GATE_4);
  not eco129 (patchNew__not_GATE_118, patchNew_new_n605_);
  nor eco130 (patchNew_new_n608_, g1015, patchNew_new_n606_);
  and eco131 (patchNew_new_n609_, patchNew__not_GATE_119, patchNew_new_n608_);
  not eco132 (patchNew__not_GATE_119, patchNew_new_n607_);
  and eco133 (patchNew_new_n611_, patchNew__not_GATE_120, g760);
  not eco134 (patchNew__not_GATE_120, g1171);
  nor eco135 (patchNew_new_n612_, patchNew_new_n289_, patchNew_new_n611_);
  and eco136 (patchNew_new_n613_, patchNew__not_GATE_121, patchNew_new_n612_);
  not eco137 (patchNew__not_GATE_121, patchNew_new_n295_);
  and eco138 (patchNew_new_n614_, g4698, patchNew_n477);
  and eco139 (patchNew_new_n615_, g839, patchNew__not_GATE_122);
  not eco140 (patchNew__not_GATE_122, patchNew_new_n613_);
  and eco141 (patchNew_new_n616_, patchNew_new_n614_, patchNew_new_n615_);
  nor eco142 (patchNew_new_n617_, patchNew_new_n401_, patchNew_new_n616_);
  nor eco143 (patchNew_new_n618_, g4795, patchNew_new_n613_);
  not eco144 (patchNew__not_GATE_21, patchNew_new_n319_);
  and eco145 (patchNew_new_n301_, g4788, g4704);
  nor eco146 (patchNew_new_n300_, g801, g730);
  nor eco147 (patchNew_new_n372_, g1015, patchNew_new_n371_);
  and eco148 (patchNew_new_n276_, g610, g608);
  not eco149 (patchNew__not_GATE_25, g730);
  and eco150 (patchNew_new_n388_, g4769, g706);
  nor eco151 (patchNew_new_n389_, patchNew_new_n385_, patchNew_new_n386_);
  and eco152 (patchNew_new_n280_, g609, g4746);
  and eco153 (patchNew_new_n341_, g625, patchNew__not_GATE_30);
  nor eco154 (patchNew_new_n438_, patchNew_new_n436_, patchNew_new_n437_);
  nor eco155 (patchNew_new_n439_, g575, patchNew_new_n364_);
  not eco156 (patchNew__not_GATE_86, patchNew_new_n461_);
  and eco157 (patchNew_new_n521_, g4802, patchNew__not_GATE_81);
  not eco158 (patchNew__not_GATE_81, patchNew_new_n519_);
  nor eco159 (patchNew_new_n522_, g509, patchNew_new_n419_);
  not eco160 (patchNew__not_GATE_33, g454);
  and eco161 (patchNew_new_n304_, g4785, patchNew__not_GATE_16);
  not eco162 (patchNew__not_GATE_15, patchNew_new_n298_);
  and eco163 (patchNew_new_n303_, patchNew_new_n301_, patchNew_new_n302_);
  and eco164 (patchNew_new_n302_, g878, g4725);
  not eco165 (patchNew__not_GATE_11, patchNew_new_n285_);
  and eco166 (patchNew_new_n286_, g753, patchNew__not_GATE_11);
  and eco167 (patchNew_new_n298_, g1024, g4736);
  nor eco168 (patchNew_new_n358_, patchNew_new_n355_, patchNew_new_n357_);
  and eco169 (patchNew_new_n299_, g625, patchNew__not_GATE_15);
  not eco170 (patchNew__not_GATE_41, patchNew_new_n373_);
  and eco171 (patchNew_new_n261_, g4721, g4754);
  not eco172 (patchNew__not_GATE_6, patchNew_new_n271_);
  not eco173 (patchNew__not_GATE_38, g4791);
  nor eco174 (patchNew_new_n348_, g4788, g1035);
  and eco175 (patchNew_new_n335_, g4785, g731);
  nor eco176 (patchNew_new_n327_, g535, patchNew_new_n326_);
  nor eco177 (patchNew_new_n285_, patchNew_new_n283_, patchNew_new_n284_);
  and eco178 (patchNew_new_n332_, g581, g4716);
  not eco179 (patchNew__not_GATE_4, patchNew_new_n266_);
  and eco180 (patchNew_new_n314_, g581, g4715);
  and eco181 (patchNew_new_n269_, g4787, patchNew__not_GATE_5);
  and eco182 (patchNew_new_n350_, g4701, patchNew_new_n309_);
  and eco183 (patchNew_new_n268_, g4815, patchNew__not_GATE_4);
  nor eco184 (patchNew_new_n349_, g4785, patchNew_new_n348_);
  nor eco185 (patchNew_new_n364_, patchNew_new_n361_, patchNew_new_n363_);
  and eco186 (patchNew_new_n322_, g804, g4738);
  not eco187 (patchNew__not_GATE_18, g4788);
  not eco188 (patchNew__not_GATE_16, patchNew_new_n303_);
  and eco189 (patchNew_new_n433_, g4680, patchNew__not_GATE_55);
  not eco190 (patchNew__not_GATE_54, patchNew_new_n431_);
  and eco191 (patchNew_new_n265_, g4732, patchNew__not_GATE_2);
  not eco192 (patchNew__not_GATE_37, patchNew_new_n361_);
  and eco193 (patchNew_new_n309_, g4785, patchNew__not_GATE_18);
  and eco194 (patchNew_new_n386_, g1122, g4749);
  not eco195 (patchNew__not_GATE_40, patchNew_new_n378_);
  and eco196 (patchNew_new_n310_, g4705, patchNew_new_n309_);
  and eco197 (patchNew_new_n313_, patchNew__not_GATE_19, patchNew_new_n312_);
  nor eco198 (patchNew_new_n380_, patchNew_new_n375_, patchNew_new_n379_);
  and eco199 (patchNew_new_n275_, g4813, patchNew__not_GATE_7);
  and eco200 (patchNew_new_n343_, g1068, g511_g4785);
  and eco201 (patchNew_new_n282_, g4813, patchNew__not_GATE_10);
  not eco202 (patchNew__not_GATE_8, patchNew_new_n273_);
  and eco203 (patchNew_new_n326_, g4785, g4707);
  and eco204 (patchNew_new_n311_, g4788, g4726);
  nor eco205 (patchNew_new_n333_, patchNew_new_n321_, patchNew_new_n332_);
  nor eco206 (patchNew_new_n281_, patchNew_new_n279_, patchNew_new_n280_);
  and eco207 (patchNew_new_n279_, g4814, g4756);
  and eco208 (patchNew_new_n356_, g4785, g4729);
  not eco209 (patchNew__not_GATE_22, patchNew_new_n322_);
  and eco210 (patchNew_new_n277_, patchNew__not_GATE_8, patchNew_new_n276_);
  and eco211 (patchNew_new_n407_, g4781, g471);
  and eco212 (patchNew_new_n330_, g542, patchNew__not_GATE_26);
  and eco213 (patchNew_new_n273_, patchNew__not_GATE_6, patchNew_new_n272_);
  not eco214 (patchNew__not_GATE_34, patchNew_new_n354_);
  and eco215 (patchNew_new_n266_, g4774, patchNew__not_GATE_3);
  nor eco216 (patchNew_new_n312_, patchNew_new_n308_, patchNew_new_n311_);
  nor eco217 (patchNew_new_n369_, g1015, patchNew_n1031);
  not eco218 (patchNew__not_GATE_0, patchNew_new_n261_);
  nor eco219 (patchNew_new_n361_, patchNew_new_n358_, patchNew_new_n360_);
  and eco220 (patchNew_new_n288_, g4814, g492);
  not eco221 (patchNew__not_GATE_31, patchNew_new_n343_);
  not eco222 (patchNew__not_GATE_32, patchNew_new_n346_);
  and eco223 (patchNew_new_n410_, g1122, g4751);
  and eco224 (patchNew_new_n319_, g4785, g4706);
  and eco225 (patchNew_new_n540_, patchNew__not_GATE_91, g4788);
  not eco226 (patchNew__not_GATE_91, g4785);
  and eco227 (patchNew_new_n541_, patchNew__not_GATE_92, g4709);
  not eco228 (patchNew__not_GATE_92, g4788);
  and eco229 (patchNew_new_n542_, g4785, patchNew__not_GATE_93);
  not eco230 (patchNew__not_GATE_93, patchNew_new_n541_);
  and eco231 (patchNew_new_n543_, g4741, g632);
  nor eco232 (patchNew_new_n544_, patchNew_new_n542_, patchNew_new_n543_);
  and eco233 (patchNew_new_n545_, g581, g4719);
  nor eco234 (patchNew_new_n546_, patchNew_new_n540_, patchNew_new_n545_);
  and eco235 (patchNew_new_n547_, patchNew__not_GATE_94, patchNew_new_n546_);
  and eco236 (patchNew_new_n548_, patchNew__not_GATE_95, patchNew_new_n547_);
  not eco237 (patchNew__not_GATE_94, patchNew_new_n544_);
  nor eco238 (patchNew_new_n429_, g510, patchNew_n1031);
  not eco239 (patchNew__not_GATE_53, patchNew_new_n427_);
  and eco240 (patchNew_new_n398_, g4773, g471);
  nor eco241 (patchNew_new_n399_, patchNew_new_n395_, patchNew_new_n396_);
  nor eco242 (patchNew_new_n400_, patchNew_new_n397_, patchNew_new_n398_);
  and eco243 (patchNew_new_n504_, patchNew_new_n502_, patchNew_new_n503_);
  and eco244 (patchNew_new_n505_, g1122, g4750);
  and eco245 (patchNew_new_n506_, g4780, g501);
  and eco246 (patchNew_new_n507_, g4770, g706);
  and eco247 (patchNew_new_n414_, patchNew__not_GATE_48, patchNew_new_n413_);
  not eco248 (patchNew__not_GATE_48, g483);
  and eco249 (patchNew_new_n492_, g4681, g460);
  and eco250 (patchNew_new_n416_, g686, patchNew_new_n415_);
  nor eco251 (patchNew_new_n345_, g1049, g1062);
  not eco252 (patchNew__not_GATE_19, patchNew_new_n310_);
  not eco253 (patchNew__not_GATE_24, patchNew_new_n327_);
  and eco254 (patchNew_new_n329_, patchNew__not_GATE_25, g4717);
  not eco255 (patchNew__not_GATE_7, patchNew_new_n274_);
  and eco256 (patchNew_new_n478_, g4775, g501);
  nor eco257 (patchNew_new_n479_, patchNew_new_n475_, patchNew_new_n476_);
  and eco258 (patchNew_new_n437_, g4799, patchNew_new_n435_);
  and eco259 (patchNew_new_n472_, patchNew__not_GATE_64, patchNew_new_n393_);
  and eco260 (patchNew_new_n468_, g4695, g483);
  not eco261 (patchNew__not_GATE_70, patchNew_new_n493_);
  not eco262 (patchNew__not_GATE_71, g4793);
  and eco263 (patchNew_new_n396_, patchNew__not_GATE_45, g4743);
  not eco264 (patchNew__not_GATE_66, g483);
  nor eco265 (patchNew_new_n483_, patchNew_new_n474_, patchNew_new_n482_);
  and eco266 (patchNew_new_n445_, g4794, patchNew__not_GATE_58);
  and eco267 (patchNew_new_n446_, g4680, patchNew_n348);
  and eco268 (patchNew_new_n424_, patchNew__not_GATE_52, patchNew_new_n423_);
  and eco269 (patchNew_new_n397_, patchNew__not_GATE_46, g706);
  not eco270 (patchNew__not_GATE_46, g555);
  nor eco271 (patchNew_new_n339_, patchNew_new_n336_, patchNew_new_n338_);
  and eco272 (patchNew_new_n283_, g4776, g705);
  and eco273 (patchNew_new_n454_, patchNew_new_n452_, patchNew_new_n453_);
  not eco274 (patchNew__not_GATE_58, patchNew_new_n441_);
  not eco275 (patchNew__not_GATE_45, g1123);
  and eco276 (patchNew_new_n354_, g576, g4740);
  nor eco277 (patchNew_new_n473_, patchNew_new_n471_, patchNew_new_n472_);
  nor eco278 (patchNew_new_n474_, g904, patchNew_new_n469_);
  and eco279 (patchNew_new_n475_, g497, g4755);
  and eco280 (patchNew_new_n336_, g730, patchNew__not_GATE_28);
  nor eco281 (patchNew_new_n305_, patchNew_new_n299_, patchNew_new_n300_);
  and eco282 (patchNew_new_n374_, g580, g4731);
  not eco283 (patchNew__not_GATE_56, g4798);
  not eco284 (patchNew__not_GATE_20, patchNew_new_n317_);
  nor eco285 (patchNew_new_n321_, patchNew_new_n318_, patchNew_new_n320_);
  and eco286 (patchNew_new_n289_, g4768, patchNew__not_GATE_12);
  nor eco287 (patchNew_new_n412_, patchNew_new_n409_, patchNew_new_n410_);
  nor eco288 (patchNew_new_n390_, patchNew_new_n387_, patchNew_new_n388_);
  and eco289 (patchNew_new_n423_, g593, patchNew__not_GATE_51);
  not eco290 (patchNew__not_GATE_49, patchNew_new_n404_);
  nor eco291 (patchNew_new_n387_, patchNew_n532, g476);
  and eco292 (patchNew_new_n462_, g685, patchNew__not_GATE_61);
  not eco293 (patchNew__not_GATE_61, patchNew_new_n415_);
  and eco294 (patchNew_new_n295_, g4813, patchNew__not_GATE_14);
  and eco295 (patchNew_new_n284_, g4814, g4766);
  and eco296 (patchNew_new_n337_, g627, g4703);
  nor eco297 (patchNew_new_n324_, patchNew_new_n316_, patchNew_new_n323_);
  and eco298 (patchNew_new_n434_, g4684, g665);
  nor eco299 (patchNew_new_n435_, patchNew_new_n433_, patchNew_new_n434_);
  not eco300 (patchNew__not_GATE_12, patchNew_new_n288_);
  not eco301 (patchNew__not_GATE_29, patchNew_new_n337_);
  and eco302 (patchNew_new_n355_, g518, patchNew__not_GATE_34);
  not eco303 (patchNew__not_GATE_10, patchNew_new_n281_);
  nor eco304 (patchNew_new_n393_, patchNew_new_n384_, patchNew_new_n392_);
  and eco305 (patchNew_new_n262_, g4711, patchNew__not_GATE_0);
  nor eco306 (patchNew_new_n448_, patchNew_new_n446_, patchNew_new_n447_);
  nor eco307 (patchNew_new_n449_, g739, patchNew_new_n448_);
  not eco308 (patchNew__not_GATE_17, patchNew_new_n304_);
  nor eco309 (patchNew_new_n365_, g4791, patchNew_new_n364_);
  not eco310 (patchNew__not_GATE_35, patchNew_new_n356_);
  and eco311 (patchNew_new_n346_, patchNew__not_GATE_31, patchNew_new_n345_);
  and eco312 (patchNew_new_n362_, g581, g4718);
  and eco313 (patchNew_new_n518_, patchNew__not_GATE_79, patchNew_n494);
  not eco314 (patchNew__not_GATE_79, g724);
  and eco315 (patchNew_new_n519_, g461, patchNew__not_GATE_80);
  not eco316 (patchNew__not_GATE_80, patchNew_new_n518_);
  and eco317 (patchNew_new_n392_, patchNew__not_GATE_43, patchNew_new_n391_);
  not eco318 (patchNew__not_GATE_43, g483);
  not eco319 (patchNew__not_GATE_13, g4814);
  and eco320 (patchNew_new_n292_, g4814, g478);
  and eco321 (patchNew_new_n290_, g4778, patchNew__not_GATE_13);
  and eco322 (patchNew_new_n421_, g569, patchNew__not_GATE_49);
  and eco323 (patchNew_new_n422_, patchNew__not_GATE_50, patchNew_n378);
  nor eco324 (patchNew_new_n480_, patchNew_new_n477_, patchNew_new_n478_);
  and eco325 (patchNew_new_n482_, patchNew__not_GATE_66, patchNew_new_n481_);
  and eco326 (patchNew_new_n444_, g4797, patchNew__not_GATE_57);
  not eco327 (patchNew__not_GATE_57, patchNew_new_n423_);
  nor eco328 (patchNew_new_n316_, g582, g730);
  not eco329 (patchNew__not_GATE_14, patchNew_new_n294_);
  not eco330 (patchNew__not_GATE_42, g4693);
  nor eco331 (patchNew_new_n382_, g4791, patchNew_n321);
  and eco332 (patchNew_new_n385_, g4779, g471);
  and eco333 (patchNew_new_n293_, g4748, g4758);
  and eco334 (patchNew_new_n484_, g4691, patchNew__not_GATE_67);
  and eco335 (patchNew_new_n485_, g4694, g600);
  not eco336 (patchNew__not_GATE_67, patchNew_n477);
  and eco337 (patchNew_new_n395_, g497, g4753);
  nor eco338 (patchNew_new_n366_, g1015, patchNew_n373);
  and eco339 (patchNew_new_n417_, g4680, patchNew_n448);
  and eco340 (patchNew_new_n418_, g4674, g460);
  not eco341 (patchNew__not_GATE_28, patchNew_new_n335_);
  and eco342 (patchNew_new_n264_, g4700, g4744);
  and eco343 (patchNew_new_n263_, g4764, patchNew__not_GATE_1);
  nor eco344 (patchNew_new_n431_, patchNew_new_n429_, patchNew_new_n430_);
  and eco345 (patchNew_new_n432_, g4798, patchNew__not_GATE_54);
  nor eco346 (patchNew_new_n352_, g448, patchNew_new_n351_);
  not eco347 (patchNew__not_GATE_3, patchNew_new_n265_);
  and eco348 (patchNew_new_n379_, g4785, patchNew__not_GATE_40);
  and eco349 (patchNew_new_n450_, patchNew__not_GATE_59, patchNew_new_n448_);
  not eco350 (patchNew__not_GATE_59, g4800);
  and eco351 (patchNew_new_n376_, g4788, g4699);
  not eco352 (patchNew__not_GATE_39, patchNew_new_n374_);
  nor eco353 (patchNew_new_n411_, patchNew_new_n407_, patchNew_new_n408_);
  nor eco354 (patchNew_new_n296_, patchNew_new_n291_, patchNew_new_n295_);
  and eco355 (patchNew_new_n340_, g630, g4735);
  not eco356 (patchNew__not_GATE_50, g533);
  and eco357 (patchNew_new_n271_, g4814, g495);
  not eco358 (patchNew__not_GATE_30, patchNew_new_n340_);
  nor eco359 (patchNew_new_n404_, patchNew_new_n402_, patchNew_new_n403_);
  nor eco360 (patchNew_new_n351_, patchNew_new_n349_, patchNew_new_n350_);
  nor eco361 (patchNew_new_n436_, g4799, patchNew_new_n435_);
  and eco362 (patchNew_new_n447_, g4685, g643);
  and eco363 (patchNew_new_n318_, g4788, patchNew__not_GATE_20);
  and eco364 (patchNew_new_n294_, patchNew_new_n292_, patchNew_new_n293_);
  and eco365 (patchNew_new_n426_, g4682, g624);
  nor eco366 (patchNew_new_n427_, patchNew_new_n425_, patchNew_new_n426_);
  nor eco367 (patchNew_new_n291_, g4813, patchNew_new_n290_);
  and eco368 (patchNew_new_n394_, g750, patchNew__not_GATE_44);
  not eco369 (patchNew__not_GATE_44, patchNew_new_n393_);
  and eco370 (patchNew_new_n363_, patchNew__not_GATE_37, patchNew_new_n362_);
  nor eco371 (patchNew_new_n307_, g4788, g648);
  not eco372 (patchNew__not_GATE_1, patchNew_new_n262_);
  xnor eco373 (patchNew__xnor_GATE_2, patchNew_new_n391_, patchNew_new_n401_);
  xnor eco374 (patchNew__xnor_GATE_3, patchNew_new_n574_, patchNew_new_n511_);
  and eco375 (patchNew_new_n451_, g550, patchNew_new_n427_);
  nor eco376 (patchNew_new_n452_, patchNew_new_n428_, patchNew_new_n449_);
  not eco377 (patchNew__not_GATE_9, patchNew_new_n275_);
  and eco378 (patchNew_new_n520_, g1332, patchNew_new_n519_);
  not eco379 (patchNew__not_GATE_64, g750);
  and eco380 (patchNew_new_n384_, patchNew__not_GATE_42, g483);
  and eco381 (patchNew_new_n368_, patchNew__not_GATE_38, patchNew_n244);
  and eco382 (patchNew_new_n317_, g4785, g4727);
  not eco383 (patchNew__not_GATE_23, patchNew_new_n321_);
  and eco384 (patchNew_new_n430_, g4683, g460);
  not eco385 (patchNew__not_GATE_51, patchNew_new_n422_);
  and eco386 (patchNew_new_n489_, g581, g4710);
  nor eco387 (patchNew_new_n490_, patchNew_new_n380_, patchNew_new_n489_);
  nor eco388 (patchNew_new_n491_, g445, patchNew_new_n490_);
  and eco389 (patchNew_new_n408_, g4771, g706);
  nor eco390 (patchNew_new_n409_, patchNew_n532, g688);
  and eco391 (patchNew_new_n420_, g509, patchNew_new_n419_);
  and eco392 (patchNew_new_n328_, g450, patchNew__not_GATE_24);
  nor eco393 (patchNew_new_n463_, g483, patchNew_n747);
  and eco394 (patchNew_new_n464_, g4689, g483);
  nor eco395 (patchNew_new_n465_, patchNew_new_n463_, patchNew_new_n464_);
  and eco396 (patchNew_new_n440_, g4672, g460);
  nor eco397 (patchNew_new_n441_, patchNew_new_n439_, patchNew_new_n440_);
  and eco398 (patchNew_new_n496_, g505, g4677);
  and eco399 (patchNew_new_n497_, patchNew__not_GATE_72, patchNew_new_n496_);
  not eco400 (patchNew__not_GATE_72, patchNew_new_n470_);
  not eco401 (patchNew__not_GATE_5, patchNew_new_n263_);
  and eco402 (patchNew_new_n359_, g536, g4708);
  not eco403 (patchNew__not_GATE_2, patchNew_new_n264_);
  and eco404 (patchNew_new_n272_, g610, g4767);
  and eco405 (patchNew_new_n510_, patchNew__not_GATE_75, patchNew_new_n509_);
  not eco406 (patchNew__not_GATE_75, patchNew_new_n508_);
  and eco407 (patchNew_new_n512_, g4691, patchNew__not_GATE_76);
  nor eco408 (patchNew_new_n419_, patchNew_new_n417_, patchNew_new_n418_);
  not eco409 (patchNew__not_GATE_55, patchNew_n770);
  and eco410 (patchNew_new_n508_, patchNew__not_GATE_74, g497);
  not eco411 (patchNew__not_GATE_74, g710);
  nor eco412 (patchNew_new_n509_, patchNew_new_n506_, patchNew_new_n507_);
  and eco413 (patchNew_new_n460_, patchNew_new_n458_, patchNew_new_n459_);
  and eco414 (patchNew_new_n461_, patchNew_new_n457_, patchNew_new_n460_);
  nor eco415 (patchNew_new_n308_, g4785, patchNew_new_n307_);
  nor eco416 (patchNew_new_n466_, g1308, patchNew_new_n465_);
  nor eco417 (patchNew_new_n467_, g553, patchNew_n1037);
  not eco418 (patchNew__not_GATE_47, g4692);
  not eco419 (patchNew__not_GATE_26, patchNew_new_n329_);
  nor eco420 (patchNew_new_n402_, g703, patchNew_new_n401_);
  and eco421 (patchNew_new_n403_, g4687, g483);
  and eco422 (patchNew_new_n360_, g4785, patchNew__not_GATE_36);
  and eco423 (patchNew_new_n274_, g4814, g4757);
  nor eco424 (patchNew_new_n373_, g633, g730);
  nor eco425 (patchNew_new_n453_, patchNew_new_n450_, patchNew_new_n451_);
  and eco426 (patchNew_new_n375_, g625, patchNew__not_GATE_39);
  and eco427 (patchNew_new_n442_, g771, patchNew_new_n441_);
  and eco428 (patchNew_new_n443_, patchNew__not_GATE_56, patchNew_new_n431_);
  and eco429 (patchNew_new_n378_, patchNew_new_n376_, patchNew_new_n377_);
  not eco430 (patchNew__not_GATE_27, patchNew_new_n330_);
  not eco431 (patchNew__not_GATE_36, patchNew_new_n359_);
  nor eco432 (patchNew_new_n469_, patchNew_new_n467_, patchNew_new_n468_);
  and eco433 (patchNew_new_n470_, patchNew__not_GATE_62, patchNew_new_n469_);
  and eco434 (patchNew_new_n428_, g4796, patchNew__not_GATE_53);
  and eco435 (patchNew_new_n338_, g4785, patchNew__not_GATE_29);
  and eco436 (patchNew_new_n323_, g625, patchNew__not_GATE_22);
  not eco437 (patchNew__not_GATE_76, patchNew_new_n511_);
  and eco438 (patchNew_new_n513_, g4688, g687);
  nor eco439 (patchNew_new_n514_, patchNew_new_n512_, patchNew_new_n513_);
  and eco440 (patchNew_new_n515_, g720, patchNew__not_GATE_77);
  not eco441 (patchNew__not_GATE_69, patchNew_new_n486_);
  not eco442 (patchNew__not_GATE_68, g4809);
  and eco443 (patchNew_new_n405_, g4803, patchNew_new_n404_);
  and eco444 (patchNew_new_n406_, patchNew__not_GATE_47, g483);
  and eco445 (patchNew_new_n457_, patchNew__not_GATE_60, patchNew_new_n456_);
  not eco446 (patchNew__not_GATE_60, patchNew_new_n444_);
  not eco447 (patchNew__not_GATE_62, g4810);
  and eco448 (patchNew_new_n471_, patchNew__not_GATE_63, patchNew_new_n465_);
  not eco449 (patchNew__not_GATE_63, g4808);
  nor eco450 (patchNew_new_n476_, g491, g1123);
  and eco451 (patchNew_new_n477_, g706, patchNew__not_GATE_65);
  not eco452 (patchNew__not_GATE_65, g487);
  and eco453 (patchNew_new_n377_, g538, g4720);
  not eco454 (patchNew__not_GATE_77, patchNew_new_n514_);
  and eco455 (patchNew_new_n516_, patchNew__not_GATE_78, patchNew_new_n514_);
  nor eco456 (patchNew_new_n517_, patchNew_new_n515_, patchNew_new_n516_);
  not eco457 (patchNew__not_GATE_78, g720);
  and eco458 (patchNew_new_n357_, g4788, patchNew__not_GATE_35);
  and eco459 (patchNew_new_n458_, patchNew_new_n454_, patchNew_new_n455_);
  nor eco460 (patchNew_new_n459_, patchNew_new_n442_, patchNew_new_n445_);
  nor eco461 (patchNew_new_n527_, patchNew_new_n421_, patchNew_new_n462_);
  and eco462 (patchNew_new_n528_, patchNew_new_n526_, patchNew_new_n527_);
  and eco463 (patchNew_new_n529_, patchNew_new_n525_, patchNew_new_n528_);
  and eco464 (patchNew_new_n530_, patchNew__not_GATE_83, patchNew_new_n529_);
  not eco465 (patchNew__not_GATE_83, patchNew_new_n517_);
  and eco466 (patchNew_new_n502_, patchNew_new_n500_, patchNew__xnor_GATE_7);
  and eco467 (patchNew_new_n503_, patchNew__not_GATE_73, patchNew_new_n499_);
  not eco468 (patchNew__not_GATE_73, patchNew_new_n473_);
  and eco469 (patchNew_new_n523_, patchNew__not_GATE_82, patchNew_new_n522_);
  not eco470 (patchNew__not_GATE_82, patchNew_new_n521_);
  nor eco471 (patchNew_new_n524_, patchNew_new_n520_, patchNew_new_n523_);
  nor eco472 (patchNew_new_n525_, patchNew_new_n394_, patchNew_new_n405_);
  nor eco473 (patchNew_new_n526_, patchNew_new_n416_, patchNew_new_n420_);
  and eco474 (patchNew_new_n425_, g4680, patchNew_n244);
  not eco475 (patchNew__not_GATE_52, g4797);
  nor eco476 (patchNew_new_n344_, g4788, g4702_g4785);
  nor eco477 (patchNew_new_n455_, patchNew_new_n424_, patchNew_new_n432_);
  nor eco478 (patchNew_new_n456_, patchNew_new_n438_, patchNew_new_n443_);
  nor eco479 (patchNew_new_n415_, patchNew_new_n406_, patchNew_new_n414_);
  and eco480 (patchNew_new_n499_, patchNew_new_n497_, patchNew__xnor_GATE_6);
  nor eco481 (patchNew_new_n500_, patchNew_new_n466_, patchNew_new_n483_);
  and eco482 (patchNew_new_n531_, patchNew__not_GATE_84, patchNew_new_n530_);
  not eco483 (patchNew__not_GATE_84, patchNew_new_n524_);
  and eco484 (patchNew_new_n532_, patchNew__not_GATE_85, patchNew_new_n531_);
  not eco485 (patchNew__not_GATE_98, patchNew_n1037);
  not eco486 (patchNew__not_GATE_85, patchNew_new_n504_);
  not eco487 (patchNew__not_GATE_95, patchNew_new_n539_);
  nor eco488 (patchNew_new_n549_, g4790, patchNew__xnor_GATE_9);
  and eco489 (patchNew_new_n550_, g864, patchNew__not_GATE_96);
  not eco490 (patchNew__not_GATE_96, patchNew_new_n547_);
  and eco491 (patchNew_new_n551_, patchNew__not_GATE_97, patchNew_new_n550_);
  not eco492 (patchNew__not_GATE_97, patchNew_new_n549_);
  not eco493 (patchNew__not_GATE_99, patchNew_n477);
  and eco494 (patchNew_new_n556_, patchNew_new_n481_, patchNew__xnor_GATE_8);
  nor eco495 (patchNew_new_n557_, patchNew_new_n481_, patchNew__xnor_GATE_8);
  nor eco496 (patchNew_new_n558_, patchNew_new_n556_, patchNew_new_n557_);
  and eco497 (patchNew_new_n534_, patchNew_new_n364_, patchNew__not_GATE_87);
  not eco498 (patchNew__not_GATE_87, patchNew_new_n490_);
  not eco499 (patchNew__not_GATE_88, patchNew_new_n371_);
  not eco500 (patchNew__not_GATE_89, patchNew_new_n535_);
  and eco501 (patchNew_new_n539_, patchNew__not_GATE_90, patchNew__xnor_GATE_9);
  not eco502 (patchNew__not_GATE_90, g4790);
  and eco503 (patchNew_new_n619_, patchNew_n477, patchNew__not_GATE_123);
  not eco504 (patchNew__not_GATE_123, patchNew_new_n618_);
  and eco505 (patchNew_new_n620_, g4698, patchNew__not_GATE_124);
  not eco506 (patchNew__not_GATE_124, patchNew_new_n619_);
  and eco507 (patchNew_new_n621_, g569, patchNew_new_n620_);
  and eco508 (patchNew_new_n622_, patchNew_new_n617_, patchNew_new_n621_);
  and eco509 (patchNew_new_n623_, patchNew_new_n413_, patchNew_new_n622_);
  and eco510 (patchNew_new_n624_, g685, patchNew__not_GATE_125);
  not eco511 (patchNew__not_GATE_125, patchNew_new_n413_);
  and eco512 (patchNew_new_n625_, patchNew__not_GATE_126, patchNew_new_n413_);
  not eco513 (patchNew__not_GATE_126, g685);
  nor eco514 (patchNew_new_n626_, patchNew_new_n624_, patchNew_new_n625_);
  and eco515 (patchNew_new_n627_, patchNew__not_GATE_127, patchNew_new_n626_);
  not eco516 (patchNew__not_GATE_127, patchNew_new_n616_);
  and eco517 (patchNew_new_n628_, patchNew_new_n620_, patchNew__not_GATE_128);
  not eco518 (patchNew__not_GATE_128, patchNew_new_n627_);
  nor eco519 (patchNew_new_n629_, patchNew_new_n623_, patchNew_new_n628_);
  and eco520 (patchNew_new_n630_, g720, patchNew__not_GATE_129);
  not eco521 (patchNew__not_GATE_129, patchNew_new_n511_);
  and eco522 (patchNew_new_n631_, patchNew__not_GATE_130, patchNew_new_n511_);
  not eco523 (patchNew__not_GATE_130, g720);
  nor eco524 (patchNew_new_n632_, patchNew_new_n630_, patchNew_new_n631_);
  and eco525 (patchNew_new_n633_, patchNew__not_GATE_131, patchNew_new_n632_);
  not eco526 (patchNew__not_GATE_131, patchNew_new_n616_);
  and eco527 (patchNew_new_n634_, patchNew_new_n620_, patchNew_new_n633_);
  and eco528 (patchNew_new_n635_, patchNew__not_GATE_132, patchNew_new_n511_);
  not eco529 (patchNew__not_GATE_132, patchNew_new_n413_);
  and eco530 (patchNew_new_n636_, patchNew_new_n620_, patchNew_new_n635_);
  and eco531 (patchNew_new_n637_, patchNew_new_n634_, patchNew__not_GATE_133);
  not eco532 (patchNew__not_GATE_133, patchNew_new_n636_);
  nor eco533 (patchNew_new_n638_, patchNew_new_n629_, patchNew_new_n637_);
  and eco534 (patchNew_new_n639_, g1332, patchNew_new_n620_);
  and eco535 (patchNew_new_n640_, patchNew__not_GATE_134, patchNew_new_n639_);
  not eco536 (patchNew__not_GATE_134, patchNew_new_n616_);
  and eco537 (patchNew_new_n641_, patchNew__not_GATE_135, patchNew_new_n640_);
  not eco538 (patchNew__not_GATE_135, patchNew_n494);
  and eco539 (patchNew_new_n642_, patchNew_new_n614_, patchNew_new_n618_);
  and eco540 (patchNew_new_n643_, g509, patchNew__not_GATE_136);
  not eco541 (patchNew__not_GATE_136, patchNew_new_n642_);
  and eco542 (patchNew_new_n644_, g4676, patchNew__not_GATE_137);
  not eco543 (patchNew__not_GATE_137, patchNew_new_n643_);
  and eco544 (patchNew_new_n645_, g4676, patchNew__not_GATE_138);
  not eco545 (patchNew__not_GATE_138, patchNew_new_n616_);
  and eco546 (patchNew_new_n646_, patchNew_n448, patchNew__not_GATE_139);
  not eco547 (patchNew__not_GATE_139, patchNew_new_n645_);
  and eco548 (patchNew_new_n647_, patchNew__not_GATE_140, patchNew_new_n646_);
  not eco549 (patchNew__not_GATE_140, patchNew_new_n644_);
  and eco550 (patchNew_new_n648_, g739, patchNew__not_GATE_141);
  not eco551 (patchNew__not_GATE_141, patchNew_new_n642_);
  and eco552 (patchNew_new_n649_, g4676, patchNew__not_GATE_142);
  not eco553 (patchNew__not_GATE_142, patchNew_new_n648_);
  and eco554 (patchNew_new_n650_, patchNew_n348, patchNew__not_GATE_143);
  not eco555 (patchNew__not_GATE_143, patchNew_new_n645_);
  and eco556 (patchNew_new_n651_, patchNew_new_n649_, patchNew__not_GATE_144);
  not eco557 (patchNew__not_GATE_144, patchNew_new_n650_);
  and eco558 (patchNew_new_n652_, g658, patchNew__not_GATE_145);
  not eco559 (patchNew__not_GATE_145, patchNew_new_n642_);
  and eco560 (patchNew_new_n653_, g618, patchNew_new_n642_);
  nor eco561 (patchNew_new_n654_, patchNew_new_n652_, patchNew_new_n653_);
  and eco562 (patchNew_new_n655_, patchNew__not_GATE_146, patchNew_new_n654_);
  not eco563 (patchNew__not_GATE_146, patchNew_n1031);
  and eco564 (patchNew_new_n656_, patchNew_n1031, patchNew__not_GATE_147);
  not eco565 (patchNew__not_GATE_147, patchNew_new_n654_);
  and eco566 (patchNew_new_n657_, g813, patchNew__not_GATE_148);
  not eco567 (patchNew__not_GATE_148, patchNew_new_n642_);
  and eco568 (patchNew_new_n658_, g790, patchNew_new_n642_);
  not eco569 (patchNew__not_GATE_149, patchNew_new_n659_);
  not eco570 (patchNew__not_GATE_150, patchNew_n770);
  nor eco571 (patchNew_new_n662_, patchNew_new_n655_, patchNew_new_n656_);
  and eco572 (patchNew_new_n664_, patchNew_new_n662_, patchNew__xnor_GATE_10);
  and eco573 (patchNew_new_n665_, patchNew_new_n651_, patchNew__not_GATE_151);
  not eco574 (patchNew__not_GATE_151, patchNew_new_n664_);
  and eco575 (patchNew_new_n666_, patchNew__not_GATE_152, patchNew_new_n650_);
  not eco576 (patchNew__not_GATE_152, patchNew_new_n649_);
  and eco577 (patchNew_new_n667_, patchNew_new_n656_, patchNew_new_n666_);
  nor eco578 (patchNew_new_n668_, patchNew_new_n665_, patchNew_new_n667_);
  and eco579 (patchNew_new_n669_, g4676, patchNew__not_GATE_153);
  not eco580 (patchNew__not_GATE_153, patchNew_new_n668_);
  and eco581 (patchNew_new_n670_, g4796, patchNew__not_GATE_154);
  not eco582 (patchNew__not_GATE_154, patchNew_new_n616_);
  and eco583 (patchNew_new_n671_, g4807, patchNew_new_n616_);
  nor eco584 (patchNew_new_n672_, patchNew_new_n670_, patchNew_new_n671_);
  and eco585 (patchNew_new_n673_, patchNew__not_GATE_155, patchNew_new_n672_);
  not eco586 (patchNew__not_GATE_155, patchNew_n244);
  and eco587 (patchNew_new_n674_, g4806, patchNew_new_n616_);
  and eco588 (patchNew_new_n675_, g4794, patchNew__not_GATE_156);
  not eco589 (patchNew__not_GATE_156, patchNew_new_n616_);
  and eco590 (patchNew_new_n676_, patchNew_n244, patchNew__not_GATE_157);
  not eco591 (patchNew__not_GATE_157, patchNew_new_n672_);
  nor eco592 (patchNew_new_n677_, patchNew_new_n674_, patchNew_new_n675_);
  and eco593 (patchNew_new_n678_, patchNew__not_GATE_158, patchNew_new_n677_);
  not eco594 (patchNew__not_GATE_158, patchNew_new_n676_);
  and eco595 (patchNew_new_n679_, patchNew_new_n364_, patchNew__not_GATE_159);
  not eco596 (patchNew__not_GATE_159, patchNew_new_n678_);
  nor eco597 (patchNew_new_n680_, patchNew_new_n673_, patchNew_new_n679_);
  and eco598 (patchNew_new_n681_, patchNew_new_n651_, patchNew__not_GATE_160);
  not eco599 (patchNew__not_GATE_160, patchNew_new_n680_);
  nor eco600 (patchNew_new_n682_, patchNew_new_n669_, patchNew_new_n681_);
  nor eco601 (patchNew_new_n683_, patchNew_new_n647_, patchNew_new_n682_);
  and eco602 (patchNew_new_n684_, patchNew__not_GATE_161, patchNew_new_n621_);
  not eco603 (patchNew__not_GATE_161, patchNew_new_n616_);
  and eco604 (patchNew_new_n685_, patchNew__not_GATE_162, patchNew_new_n620_);
  not eco605 (patchNew__not_GATE_162, patchNew_new_n617_);
  and eco606 (patchNew_new_n686_, patchNew__not_GATE_163, patchNew_new_n685_);
  not eco607 (patchNew__not_GATE_163, patchNew_new_n684_);
  nor eco608 (patchNew_new_n687_, patchNew_new_n622_, patchNew_new_n686_);
  and eco609 (patchNew_new_n688_, patchNew_new_n644_, patchNew__not_GATE_164);
  not eco610 (patchNew__not_GATE_164, patchNew_new_n646_);
  and eco611 (patchNew_new_n689_, patchNew_n494, patchNew__not_GATE_165);
  not eco612 (patchNew__not_GATE_165, patchNew_new_n616_);
  and eco613 (patchNew_new_n690_, patchNew_new_n620_, patchNew_new_n689_);
  and eco614 (patchNew_new_n691_, patchNew__not_GATE_166, patchNew_new_n690_);
  not eco615 (patchNew__not_GATE_166, patchNew_new_n639_);
  nor eco616 (patchNew_new_n692_, patchNew_new_n634_, patchNew_new_n688_);
  and eco617 (patchNew_new_n693_, patchNew__not_GATE_167, patchNew_new_n692_);
  not eco618 (patchNew__not_GATE_167, patchNew_new_n691_);
  and eco619 (patchNew_new_n694_, patchNew__not_GATE_168, patchNew_new_n693_);
  not eco620 (patchNew__not_GATE_168, patchNew_new_n641_);
  and eco621 (patchNew_new_n695_, patchNew_new_n687_, patchNew_new_n694_);
  and eco622 (patchNew_new_n696_, patchNew__not_GATE_169, patchNew_new_n695_);
  not eco623 (patchNew__not_GATE_169, patchNew_new_n683_);
  and eco624 (patchNew_new_n697_, patchNew__not_GATE_170, patchNew_new_n640_);
  not eco625 (patchNew__not_GATE_170, patchNew_new_n632_);
  nor eco626 (patchNew_new_n698_, patchNew_new_n690_, patchNew_new_n697_);
  and eco627 (patchNew_new_n699_, patchNew_new_n687_, patchNew_new_n698_);
  nor eco628 (patchNew_new_n700_, patchNew_new_n696_, patchNew_new_n699_);
  nor eco629 (patchNew_new_n701_, patchNew_new_n628_, patchNew_new_n700_);
  nor eco630 (patchNew_new_n703_, patchNew_new_n587_, patchNew_new_n591_);
  and eco631 (patchNew_new_n704_, patchNew_new_n587_, patchNew_new_n591_);
  and eco632 (patchNew_new_n706_, g581, g4715);
  and eco633 (patchNew_new_n707_, patchNew_new_n313_, patchNew__not_GATE_171);
  not eco634 (patchNew__not_GATE_171, patchNew_new_n706_);
  and eco635 (patchNew_new_n708_, patchNew__not_GATE_172, patchNew_new_n707_);
  not eco636 (patchNew__not_GATE_172, patchNew_n373);
  nor eco637 (patchNew_new_n709_, patchNew_n378, patchNew_new_n707_);
  not eco638 (patchNew__not_GATE_173, patchNew_new_n710_);
  not eco639 (patchNew__not_GATE_174, patchNew_new_n705_);
  and eco640 (patchNew_new_n714_, patchNew__not_GATE_175, patchNew__xnor_GATE_11);
  not eco641 (patchNew__not_GATE_175, patchNew_new_n605_);
  and eco642 (patchNew_new_n715_, patchNew_new_n605_, patchNew__not_GATE_176);
  not eco643 (patchNew__not_GATE_176, patchNew__xnor_GATE_11);
  nor eco644 (patchNew_new_n716_, g4697, patchNew_new_n714_);
  not eco645 (patchNew__not_GATE_177, patchNew_new_n716_);
  nor eco646 (patchNew_new_n718_, g923, g1240);
  and eco647 (patchNew_new_n719_, patchNew__not_GATE_178, patchNew_new_n718_);
  not eco648 (patchNew__not_GATE_178, patchNew_n1001);
  and eco649 (patchNew_new_n720_, g953, patchNew_n593);
  and eco650 (patchNew_new_n721_, patchNew_n835, patchNew_new_n720_);
  not eco651 (patchNew__not_GATE_179, patchNew_new_n719_);
  not eco652 (patchNew__not_GATE_180, patchNew_new_n481_);
  not eco653 (patchNew__not_GATE_181, g4811);
  not eco654 (patchNew__not_GATE_183, g4784);
  and eco655 (patchNew_new_n729_, g4669, g4671);
  and eco656 (patchNew_new_n730_, g4789, patchNew__not_GATE_182);
  not eco657 (patchNew__not_GATE_182, patchNew_new_n729_);
  and eco658 (patchNew_new_n732_, g4807, g4808);
  xnor eco659 (patchNew__xnor_GATE_0, g4811, patchNew_new_n481_);
  xnor eco660 (patchNew__xnor_GATE_1, patchNew_n747, patchNew_new_n413_);
  not eco661 (patchNew__not_GATE_184, g4809);
  and eco662 (patchNew_n477, patchNew__not_GATE_9, patchNew_new_n277_);
  nor eco663 (patchNew_n1037, patchNew_new_n282_, patchNew_new_n286_);
  nor eco664 (patchNew_n747, patchNew_new_n289_, patchNew_new_n296_);
  and eco665 (patchNew_n770, patchNew__not_GATE_17, patchNew_new_n305_);
  or eco666 (patchNew_n348, patchNew_new_n339_, patchNew_new_n341_);
  or eco667 (patchNew_n494, patchNew__not_GATE_33, patchNew_new_n352_);
  and eco668 (patchNew_new_n371_, g1340, patchNew_new_n364_);
  nor eco669 (patchNew_new_n587_, patchNew_n321, patchNew_new_n586_);
  nor eco670 (patchNew_new_n593_, patchNew_new_n588_, patchNew_new_n592_);
  nor eco671 (patchNew_new_n486_, patchNew_new_n484_, patchNew_new_n485_);
  nor eco672 (patchNew_new_n493_, patchNew_new_n491_, patchNew_new_n492_);
  nor eco673 (patchNew_new_n535_, patchNew_n321, patchNew_new_n534_);
  nor eco674 (patchNew_new_n659_, patchNew_new_n657_, patchNew_new_n658_);
  nor eco675 (patchNew_new_n705_, patchNew_new_n703_, patchNew_new_n704_);
  nor eco676 (patchNew_new_n710_, patchNew_new_n708_, patchNew_new_n709_);
  and eco677 (patchNew_new_n413_, patchNew_new_n411_, patchNew_new_n412_);
  and eco678 (patchNew_new_n391_, patchNew_new_n389_, patchNew_new_n390_);
  and eco679 (patchNew_new_n401_, patchNew_new_n399_, patchNew_new_n400_);
  nor eco680 (patchNew_new_n574_, patchNew_new_n572_, patchNew_new_n573_);
  nor eco681 (patchNew_new_n511_, patchNew_new_n505_, patchNew_new_n510_);
  nand eco682 (patchNew_n532, g4813, g4814);
  and eco683 (patchNew_new_n481_, patchNew_new_n479_, patchNew_new_n480_);
endmodule
