module top_eco(n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n21, n22, n23, n24, n25, n77, n78, n79, n80, n82, n85, n87, n98, n100, n105, n107, n108, n114, n116, n117, n119, n122, n123, n25_n23, n130, n133, n134, n135, n137, n144, n149, n152, n160_n163, n182, n189, n84_n187, n192, n23_n22, n212, n216, n218, n222, n223, n228, n233, n240, n247, n248, n253, n254, n257, n260, n267, n25_n103, n276, n288, n300, n310, n316, n317, n323, n332, n27, n28, n29, n31, n33, n35, n37, n39, n40, n42, n43, n52, n60, n64, n321, n339, n334, n336, n337, n330, n275, n314);
  input n2, n3, n4, n5;
  input n6, n7, n8, n9, n10;
  input n11, n12, n13, n14, n15;
  input n16, n17, n18, n19, n21;
  input n22, n23, n24, n25, n77;
  input n78, n79, n80, n82, n85;
  input n87, n98, n100, n105, n107;
  input n108, n114, n116, n117, n119;
  input n122, n123, n25_n23, n130, n133;
  input n134, n135, n137, n144, n149;
  input n152, n160_n163, n182, n189, n84_n187;
  input n192, n23_n22, n212, n216, n218;
  input n222, n223, n228, n233, n240;
  input n247, n248, n253, n254, n257;
  input n260, n267, n25_n103, n276, n288;
  input n300, n310, n316, n317, n323;
  input n332;
  output n27, n28, n29, n31;
  output n33, n35, n37, n39, n40;
  output n42, n43, n52, n60, n64;
  output n321, n339, n334, n336, n337;
  output n330, n275, n314;
  buf eco1 (n27, patchNew_n382);
  buf eco2 (n28, patchNew_n383);
  buf eco3 (n29, patchNew_n378);
  buf eco4 (n31, patchNew_n394);
  buf eco5 (n33, patchNew_n288);
  buf eco6 (n35, patchNew_n304);
  buf eco7 (n37, patchNew_n85);
  buf eco8 (n39, patchNew_n304);
  buf eco9 (n40, patchNew_n386);
  buf eco10 (n42, patchNew_n397);
  buf eco11 (n43, patchNew_n175);
  buf eco12 (n52, patchNew_n247);
  buf eco13 (n60, patchNew_n376);
  buf eco14 (n64, patchNew_n177);
  nand eco15 (n321, patchNew_n347, patchNew_n350);
  not eco16 (n339, patchNew_n346);
  nor eco17 (n334, patchNew_n391, patchNew_n392);
  and eco18 (n336, patchNew_n85, n11);
  not eco19 (n337, patchNew_n391);
  nor eco20 (n330, patchNew_n212_n388, n14);
  nor eco21 (n275, patchNew_n332, n16);
  nor eco22 (n314, patchNew_n308, n16);
  and eco23 (patchNew_n382, patchNew_new_n116_, patchNew_new_n117_);
  nor eco24 (patchNew_n383, n13, patchNew_new_n124_);
  nor eco25 (patchNew_n378, n130, patchNew_new_n129_);
  and eco26 (patchNew_n394, patchNew__not_GATE_9, patchNew_new_n131_);
  and eco27 (patchNew_n288, patchNew__not_GATE_12, patchNew_new_n134_);
  nor eco28 (patchNew_n304, n22, patchNew_new_n127_);
  nor eco29 (patchNew_n85, n23_n22, n135);
  and eco30 (patchNew_n386, n10, patchNew_n397);
  and eco31 (patchNew_n397, patchNew_new_n137_, patchNew_new_n138_);
  nor eco32 (patchNew_n175, n23, patchNew_new_n141_);
  nor eco33 (patchNew_n247, n16, patchNew_new_n178_);
  nor eco34 (patchNew_n376, n16, patchNew_new_n198_);
  or eco35 (patchNew_n177, patchNew_new_n206_, patchNew_new_n244_);
  and eco36 (patchNew_n308, patchNew_new_n273_, patchNew_new_n275_);
  and eco37 (patchNew_n332, patchNew__not_GATE_83, patchNew_new_n292_);
  and eco38 (patchNew_n346, patchNew_new_n296_, patchNew_new_n297_);
  or eco39 (patchNew_n347, n152, patchNew_n346);
  nor eco40 (patchNew_n350, patchNew_new_n149_, patchNew_new_n300_);
  and eco41 (patchNew_n212_n388, n130, patchNew_new_n302_);
  nand eco42 (patchNew_n391, n119, patchNew_new_n137_);
  nand eco43 (patchNew_n392, n14, n21);
  nor eco44 (patchNew_new_n173_, patchNew_new_n170_, patchNew_new_n172_);
  nor eco45 (patchNew_new_n174_, n134, patchNew_n386);
  and eco46 (patchNew_new_n175_, patchNew__not_GATE_26, patchNew_new_n174_);
  not eco47 (patchNew__not_GATE_26, patchNew_new_n173_);
  and eco48 (patchNew_new_n121_, n9, patchNew__not_GATE_6);
  and eco49 (patchNew_new_n127_, patchNew__not_GATE_8, patchNew_new_n126_);
  nor eco50 (patchNew_new_n115_, n107, patchNew_new_n110_);
  and eco51 (patchNew_new_n120_, n7, patchNew__not_GATE_5);
  not eco52 (patchNew__not_GATE_3, patchNew_new_n112_);
  and eco53 (patchNew_new_n143_, n134, n25);
  not eco54 (patchNew__not_GATE_14, patchNew_new_n148_);
  not eco55 (patchNew__not_GATE_10, n11);
  not eco56 (patchNew__not_GATE_2, n23);
  and eco57 (patchNew_new_n133_, patchNew__not_GATE_10, n21);
  not eco58 (patchNew__not_GATE_6, patchNew_new_n120_);
  not eco59 (patchNew__not_GATE_24, n19);
  and eco60 (patchNew_new_n172_, patchNew__not_GATE_25, patchNew_new_n171_);
  not eco61 (patchNew__not_GATE_25, n25);
  and eco62 (patchNew_new_n162_, n23, patchNew__not_GATE_21);
  not eco63 (patchNew__not_GATE_21, patchNew_new_n161_);
  not eco64 (patchNew__not_GATE_4, patchNew_new_n114_);
  and eco65 (patchNew_new_n131_, n134, n21);
  and eco66 (patchNew_new_n116_, patchNew__not_GATE_4, patchNew_new_n115_);
  and eco67 (patchNew_new_n112_, n22, patchNew_new_n111_);
  and eco68 (patchNew_new_n152_, n218, patchNew__not_GATE_16);
  not eco69 (patchNew__not_GATE_7, patchNew_n224);
  and eco70 (patchNew_new_n117_, n323, n117);
  not eco71 (patchNew__not_GATE_5, patchNew_new_n119_);
  and eco72 (patchNew_new_n111_, n12, patchNew__not_GATE_1);
  and eco73 (patchNew_new_n134_, n22, patchNew__not_GATE_11);
  and eco74 (patchNew_new_n114_, patchNew__not_GATE_3, patchNew_new_n113_);
  and eco75 (patchNew_new_n150_, patchNew__not_GATE_15, patchNew_new_n124_);
  and eco76 (patchNew_new_n151_, n108, n133);
  and eco77 (patchNew_new_n113_, patchNew__not_GATE_2, n218);
  not eco78 (patchNew__not_GATE_12, patchNew_new_n133_);
  nor eco79 (patchNew_new_n129_, n123, patchNew_n304);
  and eco80 (patchNew_new_n110_, n228, patchNew__not_GATE_0);
  not eco81 (patchNew__not_GATE_9, n260);
  not eco82 (patchNew__not_GATE_8, n332);
  nor eco83 (patchNew_new_n165_, patchNew_new_n155_, patchNew_new_n164_);
  nor eco84 (patchNew_new_n161_, n253, patchNew_new_n160_);
  and eco85 (patchNew_new_n119_, n2, n3);
  and eco86 (patchNew_new_n126_, n23, n24);
  not eco87 (patchNew__not_GATE_23, patchNew_new_n167_);
  nor eco88 (patchNew_new_n170_, n13, n135);
  and eco89 (patchNew_new_n171_, patchNew__not_GATE_24, patchNew_n210);
  and eco90 (patchNew_new_n144_, n160_n163, patchNew_new_n143_);
  nor eco91 (patchNew_new_n155_, n189, patchNew_new_n154_);
  not eco92 (patchNew__not_GATE_15, n13);
  and eco93 (patchNew_new_n160_, n78, patchNew_new_n159_);
  not eco94 (patchNew__not_GATE_18, n7);
  not eco95 (patchNew__not_GATE_13, n79);
  and eco96 (patchNew_new_n122_, patchNew__not_GATE_7, patchNew_new_n121_);
  nor eco97 (patchNew_new_n156_, n87, patchNew_new_n137_);
  and eco98 (patchNew_new_n157_, n144, patchNew__not_GATE_18);
  and eco99 (patchNew_new_n158_, n3, patchNew__not_GATE_19);
  nor eco100 (patchNew_new_n137_, n23, n24);
  not eco101 (patchNew__not_GATE_0, n6);
  nor eco102 (patchNew_new_n123_, n310, patchNew_new_n122_);
  not eco103 (patchNew__not_GATE_1, n21);
  and eco104 (patchNew_new_n149_, patchNew_new_n145_, patchNew__not_GATE_14);
  not eco105 (patchNew__not_GATE_11, n25_n23);
  not eco106 (patchNew__not_GATE_19, patchNew_new_n157_);
  and eco107 (patchNew_new_n159_, n9, patchNew__not_GATE_20);
  not eco108 (patchNew__not_GATE_20, patchNew_new_n158_);
  nor eco109 (patchNew_new_n192_, n182, n17);
  not eco110 (patchNew__not_GATE_27, patchNew_new_n169_);
  nor eco111 (patchNew_new_n177_, patchNew_new_n144_, patchNew_new_n149_);
  and eco112 (patchNew_new_n178_, patchNew__not_GATE_28, patchNew_new_n177_);
  not eco113 (patchNew__not_GATE_28, patchNew_new_n176_);
  nor eco114 (patchNew_new_n124_, n233, patchNew_new_n123_);
  and eco115 (patchNew_new_n154_, n12, patchNew__not_GATE_17);
  not eco116 (patchNew__not_GATE_17, patchNew_new_n153_);
  nor eco117 (patchNew_new_n147_, n21, n22);
  and eco118 (patchNew_new_n148_, patchNew_new_n146_, patchNew_new_n147_);
  and eco119 (patchNew_new_n180_, patchNew__not_GATE_29, n84_n187);
  not eco120 (patchNew__not_GATE_29, n189);
  and eco121 (patchNew_new_n181_, n216, n8);
  and eco122 (patchNew_new_n182_, n218, patchNew__not_GATE_30);
  not eco123 (patchNew__not_GATE_30, patchNew_new_n181_);
  and eco124 (patchNew_new_n183_, patchNew__not_GATE_31, patchNew_new_n121_);
  not eco125 (patchNew__not_GATE_31, n192);
  nor eco126 (patchNew_new_n138_, n253, n135);
  and eco127 (patchNew_new_n176_, patchNew__not_GATE_27, patchNew_new_n175_);
  nor eco128 (patchNew_new_n166_, patchNew_new_n152_, patchNew_new_n165_);
  and eco129 (patchNew_new_n153_, n80, n79);
  not eco130 (patchNew__not_GATE_16, patchNew_new_n151_);
  nor eco131 (patchNew_new_n163_, patchNew_new_n131_, patchNew_new_n156_);
  and eco132 (patchNew_new_n164_, patchNew__not_GATE_22, patchNew_new_n163_);
  not eco133 (patchNew__not_GATE_22, patchNew_new_n162_);
  nor eco134 (patchNew_new_n145_, n24, n25);
  nor eco135 (patchNew_new_n146_, n149, n18);
  nor eco136 (patchNew_new_n167_, n116, patchNew_new_n166_);
  nor eco137 (patchNew_new_n168_, patchNew_n378, patchNew_new_n150_);
  and eco138 (patchNew_new_n169_, patchNew__not_GATE_23, patchNew_new_n168_);
  and eco139 (patchNew_new_n141_, patchNew_n173, patchNew__not_GATE_13);
  nor eco140 (patchNew_new_n184_, n233, patchNew_new_n183_);
  nor eco141 (patchNew_new_n185_, n12, n23_n22);
  and eco142 (patchNew_new_n186_, n24, patchNew_new_n185_);
  and eco143 (patchNew_new_n187_, patchNew_n360, patchNew__not_GATE_32);
  not eco144 (patchNew__not_GATE_32, patchNew_new_n186_);
  nor eco145 (patchNew_new_n188_, patchNew_new_n180_, patchNew_new_n182_);
  and eco146 (patchNew_new_n189_, patchNew__not_GATE_33, patchNew_new_n188_);
  not eco147 (patchNew__not_GATE_33, patchNew_new_n187_);
  and eco148 (patchNew_new_n190_, patchNew__not_GATE_34, patchNew_new_n189_);
  not eco149 (patchNew__not_GATE_34, patchNew_new_n184_);
  nor eco150 (patchNew_new_n191_, n116, patchNew_new_n190_);
  and eco151 (patchNew_new_n194_, n24, n137);
  and eco152 (patchNew_new_n193_, patchNew_n304, patchNew_new_n192_);
  nor eco153 (patchNew_new_n217_, n182, n16);
  and eco154 (patchNew_new_n195_, patchNew_new_n143_, patchNew_new_n194_);
  nor eco155 (patchNew_new_n196_, patchNew_n288, patchNew_new_n195_);
  and eco156 (patchNew_new_n197_, patchNew__not_GATE_35, patchNew_new_n196_);
  not eco157 (patchNew__not_GATE_35, patchNew_new_n193_);
  and eco158 (patchNew_new_n198_, patchNew__not_GATE_36, patchNew_new_n197_);
  not eco159 (patchNew__not_GATE_36, patchNew_new_n191_);
  and eco160 (patchNew_new_n200_, n10, patchNew__not_GATE_37);
  not eco161 (patchNew__not_GATE_37, n24);
  nor eco162 (patchNew_new_n201_, n23, patchNew_new_n200_);
  and eco163 (patchNew_new_n202_, n254, patchNew__not_GATE_38);
  not eco164 (patchNew__not_GATE_38, patchNew_new_n201_);
  nor eco165 (patchNew_new_n203_, n119, n248);
  and eco166 (patchNew_new_n204_, patchNew__not_GATE_39, patchNew_new_n203_);
  not eco167 (patchNew__not_GATE_39, patchNew_new_n202_);
  nor eco168 (patchNew_new_n205_, n16, patchNew_new_n204_);
  and eco169 (patchNew_new_n206_, patchNew_n175, patchNew__not_GATE_40);
  not eco170 (patchNew__not_GATE_40, patchNew_new_n205_);
  and eco171 (patchNew_new_n207_, patchNew__not_GATE_41, patchNew_new_n144_);
  not eco172 (patchNew__not_GATE_41, n16);
  and eco173 (patchNew_new_n208_, n85, patchNew_new_n145_);
  and eco174 (patchNew_new_n209_, n21, patchNew__not_GATE_42);
  not eco175 (patchNew__not_GATE_42, patchNew_new_n208_);
  and eco176 (patchNew_new_n210_, n114, patchNew_new_n209_);
  nor eco177 (patchNew_new_n211_, patchNew_n85, patchNew_new_n210_);
  nor eco178 (patchNew_new_n212_, n16, patchNew_new_n211_);
  and eco179 (patchNew_new_n213_, n82, n77);
  and eco180 (patchNew_new_n214_, n17, patchNew__not_GATE_43);
  not eco181 (patchNew__not_GATE_43, patchNew_new_n213_);
  and eco182 (patchNew_new_n215_, n25_n23, patchNew__not_GATE_44);
  not eco183 (patchNew__not_GATE_44, patchNew_new_n214_);
  and eco184 (patchNew_new_n216_, n105, patchNew__not_GATE_45);
  not eco185 (patchNew__not_GATE_45, patchNew_new_n215_);
  and eco186 (patchNew_new_n219_, patchNew__not_GATE_46, patchNew_new_n218_);
  nor eco187 (patchNew_new_n218_, n22, patchNew_new_n217_);
  and eco188 (patchNew_new_n248_, n14, patchNew__not_GATE_61);
  not eco189 (patchNew__not_GATE_46, patchNew_new_n216_);
  and eco190 (patchNew_new_n220_, n79, patchNew__not_GATE_47);
  not eco191 (patchNew__not_GATE_47, patchNew_new_n219_);
  nor eco192 (patchNew_new_n221_, patchNew_new_n212_, patchNew_new_n220_);
  and eco193 (patchNew_new_n222_, patchNew__not_GATE_48, patchNew_new_n146_);
  not eco194 (patchNew__not_GATE_48, n16);
  and eco195 (patchNew_new_n223_, patchNew_new_n147_, patchNew__not_GATE_49);
  not eco196 (patchNew__not_GATE_49, patchNew_new_n222_);
  and eco197 (patchNew_new_n224_, patchNew_new_n145_, patchNew__not_GATE_50);
  not eco198 (patchNew__not_GATE_50, patchNew_new_n223_);
  nor eco199 (patchNew_new_n225_, n13, n16);
  and eco200 (patchNew_new_n226_, n257, n114);
  and eco201 (patchNew_new_n227_, n222, n223);
  and eco202 (patchNew_new_n228_, patchNew_n125, patchNew__not_GATE_51);
  not eco203 (patchNew__not_GATE_51, patchNew_new_n227_);
  nor eco204 (patchNew_new_n229_, n212, n14);
  nor eco205 (patchNew_new_n230_, patchNew_n135, patchNew_new_n229_);
  and eco206 (patchNew_new_n231_, patchNew__not_GATE_52, patchNew_new_n230_);
  not eco207 (patchNew__not_GATE_52, patchNew_new_n228_);
  nor eco208 (patchNew_new_n232_, n100, patchNew_new_n126_);
  and eco209 (patchNew_new_n233_, n25, patchNew__not_GATE_53);
  not eco210 (patchNew__not_GATE_53, patchNew_new_n137_);
  and eco211 (patchNew_new_n234_, patchNew__not_GATE_54, patchNew_new_n233_);
  not eco212 (patchNew__not_GATE_54, patchNew_new_n232_);
  nor eco213 (patchNew_new_n235_, patchNew_new_n226_, patchNew_new_n231_);
  and eco214 (patchNew_new_n236_, patchNew__not_GATE_55, patchNew_new_n235_);
  not eco215 (patchNew__not_GATE_55, patchNew_new_n234_);
  and eco216 (patchNew_new_n237_, patchNew__not_GATE_56, patchNew_new_n236_);
  not eco217 (patchNew__not_GATE_56, patchNew_new_n116_);
  and eco218 (patchNew_new_n238_, patchNew_new_n225_, patchNew__not_GATE_57);
  not eco219 (patchNew__not_GATE_57, patchNew_new_n237_);
  nor eco220 (patchNew_new_n239_, patchNew_new_n221_, patchNew_new_n224_);
  and eco221 (patchNew_new_n240_, patchNew__not_GATE_58, patchNew_new_n239_);
  not eco222 (patchNew__not_GATE_58, patchNew_new_n238_);
  and eco223 (patchNew_new_n241_, n25, patchNew_new_n185_);
  and eco224 (patchNew_new_n242_, patchNew_new_n225_, patchNew_new_n241_);
  nor eco225 (patchNew_new_n243_, patchNew_new_n207_, patchNew_new_n242_);
  and eco226 (patchNew_new_n244_, patchNew__not_GATE_59, patchNew_new_n243_);
  not eco227 (patchNew__not_GATE_59, patchNew_new_n240_);
  and eco228 (patchNew_new_n246_, n13, patchNew__not_GATE_60);
  not eco229 (patchNew__not_GATE_60, n233);
  nor eco230 (patchNew_new_n247_, n288, patchNew_new_n209_);
  and eco231 (patchNew_new_n266_, n21, n134);
  not eco232 (patchNew__not_GATE_61, patchNew_new_n247_);
  and eco233 (patchNew_new_n249_, n310, patchNew_new_n143_);
  and eco234 (patchNew_new_n250_, patchNew__not_GATE_62, n310);
  not eco235 (patchNew__not_GATE_62, n233);
  nor eco236 (patchNew_new_n251_, n189, n152);
  and eco237 (patchNew_new_n252_, n276, patchNew_new_n131_);
  and eco238 (patchNew_new_n253_, n14, patchNew__not_GATE_63);
  not eco239 (patchNew__not_GATE_63, patchNew_new_n252_);
  and eco240 (patchNew_new_n254_, patchNew__not_GATE_64, n23);
  not eco241 (patchNew__not_GATE_64, n152);
  nor eco242 (patchNew_new_n255_, n24, n25_n103);
  and eco243 (patchNew_new_n256_, patchNew__not_GATE_65, patchNew_new_n255_);
  not eco244 (patchNew__not_GATE_65, patchNew_new_n254_);
  nor eco245 (patchNew_new_n257_, patchNew_new_n251_, patchNew_new_n256_);
  and eco246 (patchNew_new_n258_, patchNew__not_GATE_66, patchNew_new_n257_);
  not eco247 (patchNew__not_GATE_66, patchNew_new_n253_);
  nor eco248 (patchNew_new_n259_, patchNew_new_n250_, patchNew_new_n258_);
  and eco249 (patchNew_new_n260_, n4, n5);
  nor eco250 (patchNew_new_n261_, n6, patchNew_new_n260_);
  and eco251 (patchNew_new_n262_, n14, patchNew__not_GATE_67);
  not eco252 (patchNew__not_GATE_67, patchNew_new_n261_);
  and eco253 (patchNew_new_n263_, n12, patchNew_new_n152_);
  and eco254 (patchNew_new_n264_, patchNew__not_GATE_68, patchNew_new_n263_);
  not eco255 (patchNew__not_GATE_68, patchNew_new_n262_);
  nor eco256 (patchNew_new_n265_, patchNew_n397, patchNew_new_n264_);
  and eco257 (patchNew_new_n300_, n114, patchNew__not_GATE_87);
  and eco258 (patchNew_new_n267_, patchNew__not_GATE_69, n316);
  not eco259 (patchNew__not_GATE_69, n25);
  nor eco260 (patchNew_new_n268_, patchNew_new_n266_, patchNew_new_n267_);
  nor eco261 (patchNew_new_n269_, n152, patchNew_new_n268_);
  nor eco262 (patchNew_new_n270_, patchNew_n288, patchNew_new_n246_);
  and eco263 (patchNew_new_n271_, patchNew__not_GATE_70, patchNew_new_n270_);
  not eco264 (patchNew__not_GATE_70, patchNew_new_n249_);
  and eco265 (patchNew_new_n272_, patchNew__not_GATE_71, patchNew_new_n271_);
  not eco266 (patchNew__not_GATE_71, patchNew_new_n269_);
  and eco267 (patchNew_new_n273_, patchNew__not_GATE_72, patchNew_new_n272_);
  not eco268 (patchNew__not_GATE_72, patchNew_new_n193_);
  nor eco269 (patchNew_new_n274_, patchNew_new_n248_, patchNew_new_n259_);
  and eco270 (patchNew_new_n275_, patchNew__not_GATE_73, patchNew_new_n274_);
  not eco271 (patchNew__not_GATE_73, patchNew_new_n265_);
  and eco272 (patchNew_new_n277_, n257, n116);
  and eco273 (patchNew_new_n278_, n23, patchNew__not_GATE_74);
  not eco274 (patchNew__not_GATE_74, n24);
  and eco275 (patchNew_new_n279_, n100, patchNew__not_GATE_75);
  not eco276 (patchNew__not_GATE_75, patchNew_new_n159_);
  nor eco277 (patchNew_new_n280_, n116, n276);
  and eco278 (patchNew_new_n281_, patchNew__not_GATE_76, patchNew_new_n280_);
  not eco279 (patchNew__not_GATE_76, patchNew_new_n279_);
  and eco280 (patchNew_new_n282_, patchNew_new_n278_, patchNew__not_GATE_77);
  not eco281 (patchNew__not_GATE_77, patchNew_new_n281_);
  and eco282 (patchNew_new_n283_, n21, patchNew__not_GATE_78);
  not eco283 (patchNew__not_GATE_78, patchNew_new_n204_);
  and eco284 (patchNew_new_n284_, n24, patchNew_new_n192_);
  and eco285 (patchNew_new_n285_, n21, patchNew__not_GATE_79);
  not eco286 (patchNew__not_GATE_79, patchNew_new_n284_);
  nor eco287 (patchNew_new_n286_, n25_n103, patchNew_new_n285_);
  and eco288 (patchNew_new_n287_, n240, n267);
  and eco289 (patchNew_new_n288_, n189, patchNew__not_GATE_80);
  not eco290 (patchNew__not_GATE_80, patchNew_new_n287_);
  nor eco291 (patchNew_new_n289_, patchNew_n298, patchNew_new_n288_);
  nor eco292 (patchNew_new_n290_, patchNew_new_n277_, patchNew_new_n289_);
  and eco293 (patchNew_new_n291_, patchNew__not_GATE_81, patchNew_new_n290_);
  not eco294 (patchNew__not_GATE_81, patchNew_new_n286_);
  and eco295 (patchNew_new_n292_, patchNew__not_GATE_82, patchNew_new_n291_);
  not eco296 (patchNew__not_GATE_82, patchNew_new_n283_);
  not eco297 (patchNew__not_GATE_83, patchNew_new_n282_);
  and eco298 (patchNew_new_n294_, patchNew__not_GATE_84, patchNew_new_n278_);
  not eco299 (patchNew__not_GATE_84, n25_n103);
  and eco300 (patchNew_new_n295_, n189, n317);
  and eco301 (patchNew_new_n296_, patchNew__not_GATE_85, patchNew_new_n295_);
  not eco302 (patchNew__not_GATE_85, patchNew_new_n294_);
  and eco303 (patchNew_new_n297_, n233, patchNew__not_GATE_86);
  not eco304 (patchNew__not_GATE_86, patchNew_new_n266_);
  not eco305 (patchNew__not_GATE_87, patchNew_new_n296_);
  and eco306 (patchNew_new_n302_, n15, patchNew__not_GATE_88);
  not eco307 (patchNew__not_GATE_88, n122);
  nand eco308 (patchNew_n224, n12, n25);
  nor eco309 (patchNew_n210, n21, n24);
  nor eco310 (patchNew_n173, patchNew_n172, n22);
  nand eco311 (patchNew_n360, n300, patchNew_n125);
  nor eco312 (patchNew_n125, n98, n260);
  nor eco313 (patchNew_n135, n247, n212);
  nand eco314 (patchNew_n298, n12, n24);
  not eco315 (patchNew_n172, n21);
endmodule
