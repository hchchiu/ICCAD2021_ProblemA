module top_eco(\y[7]_in, \a[0], n_490, \op[0], \a[1], \a[2], \a[3], \a[4], \a[5], \b[0], \b[1], \b[2], \b[3], \b[4], \b[5], \op[1], n_505, n_506, wc1, n_474, wc3, n_482, n_489, wc7, n_534, n_535, n_549, n_544, n_569, n_573, n_665, wc52, n_713, n_698, n_668, wc37, n_683, wc42, n_472, wc47, n_471, n_710, n_582, n_725, n_680, n_695, wc61, overflow, greater, is_eq, \y[0], parity, \y[1], \y[2], \y[3], \y[4], \y[5], \y[6], \y[7], less);
  input \y[7]_in, \a[0], n_490, \op[0], \a[1];
  input \a[2], \a[3], \a[4], \a[5], \b[0];
  input \b[1], \b[2], \b[3], \b[4], \b[5];
  input \op[1], n_505, n_506, wc1, n_474;
  input wc3, n_482, n_489, wc7, n_534;
  input n_535, n_549, n_544, n_569, n_573;
  input n_665, wc52, n_713, n_698, n_668;
  input wc37, n_683, wc42, n_472, wc47;
  input n_471, n_710, n_582, n_725, n_680;
  input n_695, wc61;
  output overflow, greater, is_eq, \y[0], parity;
  output \y[1], \y[2], \y[3], \y[4], \y[5];
  output \y[6], \y[7], less;
  wire nn_539, nwc11, nn_264, nn_475, nn_496;
  wire nn_535, nn_803, nn_540, nn_541, nn_802;
  wire nwc10, nn_195, nn_451, nn_732, nwc28;
  wire nn_551, nn_804, nwc12, nn_450, nn_502;
  wire nn_805, nwc13, nn_806, nwc14, nn_193;
  wire nn_190, nn_807, nwc15, nn_536, nwc16;
  wire nn_729, nn_728, nn_714, nn_811, nn_140;
  wire nn_544, nwc29, nwc17, nn_191, nn_503;
  wire nn_812, nwc18, nn_726, nn_727, nn_69;
  wire nn_505, nwc19, nn_783, nn_782, nwc20;
  wire nwc21, nn_545, nn_711, nn_710, nwc22;
  wire nn_696, nwc23, nn_780, nn_339, nwc24;
  wire nn_701, nn_702, nn_445, nn_550, nn_455;
  wire nn_705, nn_819, nwc25, nn_194, nn_192;
  wire nn_820, nwc26, nn_694, nn_695, nn_413;
  wire nn_654, nn_185, nn_453, nn_670, nn_771;
  wire nn_770, nwc30, nwc31, nn_672, nwc32;
  wire nn_522, nn_671, nn_641, nn_687, nn_653;
  wire nwc33, nn_546, nn_683, nn_768, nn_677;
  wire nn_678, nn_47, nwc34, nn_759, nn_758;
  wire nn_636, nwc35, nwc36, nn_547, nwc37;
  wire nn_369, nwc38, nn_652, nwc39, nn_410;
  wire nn_642, nn_756, nn_634, nn_635, nn_143;
  wire nn_552, nwc40, nn_524, nn_651, nn_657;
  wire nn_662, nn_597, nwc41, nwc42, nn_553;
  wire nn_56, nn_611, nwc43, nn_747, nn_746;
  wire nn_538, nn_627, nwc44, nn_555, nwc45;
  wire nn_620, nn_602, nn_603, nn_744, nn_626;
  wire nwc46, nn_595, nn_596, nn_521, nn_615;
  wire nn_606, nn_548, nn_570, nwc47, nn_41;
  wire nn_612, nn_537, nwc48, nn_360, nwc49;
  wire nwc50, nn_549, nn_554, nn_543, nn_579;
  wire nwc51, nn_588, nn_735, nn_584, nn_575;
  wire nn_576, nn_568, nn_569, nn_561, nwc52;
  wire nwc53, nwc54, nwc55, nwc63, nwc64;
  wire nwc65, nwc66, nwc67, nwc68, nwc69;
  assign overflow = \y[7]_in;
  and eco2 (greater, nn_538, nn_339);
  and eco3 (is_eq, nn_505, nwc64);
  or eco4 (nn_539, \a[2], \b[2]);
  and eco5 (\y[0], nn_195, nwc66);
  nand eco6 (parity, nn_802, nn_803);
  and eco7 (\y[1], nn_194, nwc63);
  and eco8 (\y[2], nn_193, nwc68);
  and eco9 (\y[3], nn_192, nwc67);
  and eco10 (\y[4], nn_191, nwc65);
  and eco11 (\y[5], nwc69, nn_190);
  assign \y[6] = \y[7]_in;
  not eco13 (\y[7], nn_69);
  nand eco14 (less, n_544, nn_732);
  not eco15 (nwc11, nn_195);
  or eco16 (nn_264, wc52, \op[1]);
  or eco17 (nn_475, wc61, \a[5]);
  or eco18 (nn_496, wc42, \a[0]);
  or eco19 (nn_535, \a[4], \b[4]);
  or eco20 (nn_803, nn_451, nwc11);
  or eco21 (nn_540, \a[3], \b[3]);
  or eco22 (nn_541, \a[1], \b[1]);
  or eco23 (nn_802, nwc10, nn_195);
  not eco24 (nwc10, nn_451);
  nand eco25 (nn_195, nn_611, nn_612);
  nand eco26 (nn_451, nn_804, nn_805);
  nand eco27 (nn_732, nn_536, n_549);
  not eco28 (nwc28, nn_551);
  nand eco29 (nn_551, nn_677, nn_678);
  or eco30 (nn_804, nwc12, nn_450);
  not eco31 (nwc12, nn_502);
  nand eco32 (nn_450, nn_811, nn_812);
  nand eco33 (nn_502, nn_806, nn_807);
  or eco34 (nn_805, nn_502, nwc13);
  not eco35 (nwc13, nn_450);
  or eco36 (nn_806, nwc14, nn_193);
  not eco37 (nwc14, nn_190);
  or eco38 (nn_193, nwc34, nn_759);
  or eco39 (nn_190, nwc16, nn_729);
  or eco40 (nn_807, nn_190, nwc15);
  not eco41 (nwc15, nn_193);
  nand eco42 (nn_536, n_535, nn_714);
  not eco43 (nwc16, nn_728);
  nand eco44 (nn_729, nn_726, nn_727);
  nand eco45 (nn_728, nn_140, nn_544);
  or eco46 (nn_714, nwc20, nn_505);
  or eco47 (nn_811, nwc17, nn_191);
  nand eco48 (nn_140, nn_455, nn_475);
  or eco49 (nn_544, nn_696, nwc23);
  not eco50 (nwc29, nn_770);
  not eco51 (nwc17, nn_503);
  or eco52 (nn_191, nwc19, nn_783);
  nand eco53 (nn_503, nn_819, nn_820);
  or eco54 (nn_812, nn_503, nwc18);
  not eco55 (nwc18, nn_191);
  or eco56 (nn_726, nwc21, nn_140);
  or eco57 (nn_727, n_725, n_471);
  or eco58 (nn_69, nn_505, nn_264);
  nand eco59 (nn_505, nn_455, nn_705);
  not eco60 (nwc19, nn_782);
  nand eco61 (nn_783, nn_780, n_713);
  nand eco62 (nn_782, nn_445, nn_550);
  not eco63 (nwc20, n_534);
  not eco64 (nwc21, nn_545);
  nand eco65 (nn_545, nn_701, nn_702);
  or eco66 (nn_711, nn_710, nwc22);
  or eco67 (nn_710, nn_339, nwc24);
  not eco68 (nwc22, n_544);
  nand eco69 (nn_696, nn_694, nn_695);
  not eco70 (nwc23, n_472);
  or eco71 (nn_780, nwc28, nn_445);
  or eco72 (nn_339, nn_654, wc37);
  not eco73 (nwc24, n_535);
  or eco74 (nn_701, nn_185, nwc31);
  or eco75 (nn_702, nn_264, nn_413);
  nand eco76 (nn_445, n_482, nn_522);
  or eco77 (nn_550, nn_672, nwc32);
  or eco78 (nn_455, wc7, \b[5]);
  nand eco79 (nn_705, nn_475, nn_413);
  or eco80 (nn_819, nwc25, nn_194);
  not eco81 (nwc25, nn_192);
  or eco82 (nn_194, nwc43, nn_747);
  or eco83 (nn_192, nwc29, nn_771);
  or eco84 (nn_820, nn_192, nwc26);
  not eco85 (nwc26, nn_194);
  or eco86 (nn_694, nn_185, nn_453);
  or eco87 (nn_695, nn_264, nwc30);
  nand eco88 (nn_413, nn_522, nn_687);
  or eco89 (nn_654, nn_653, nwc33);
  or eco90 (nn_185, \op[1], \op[0]);
  nand eco91 (nn_453, nn_683, n_710);
  or eco92 (nn_670, nn_264, nwc37);
  nand eco93 (nn_771, nn_768, n_698);
  nand eco94 (nn_770, n_569, nn_546);
  not eco95 (nwc30, nn_413);
  not eco96 (nwc31, nn_453);
  nand eco97 (nn_672, nn_670, nn_671);
  not eco98 (nwc32, n_472);
  or eco99 (nn_522, wc3, \b[4]);
  or eco100 (nn_671, nn_185, nn_47);
  or eco101 (nn_641, nn_185, nwc44);
  nand eco102 (nn_687, n_482, nn_369);
  or eco103 (nn_653, nn_652, nwc39);
  not eco104 (nwc33, nn_522);
  or eco105 (nn_546, nn_636, nwc35);
  nand eco106 (nn_683, nn_535, nn_47);
  or eco107 (nn_768, nwc36, n_569);
  or eco108 (nn_677, nn_185, nwc38);
  or eco109 (nn_678, nn_264, nn_369);
  nand eco110 (nn_47, nn_662, n_695);
  not eco111 (nwc34, nn_758);
  nand eco112 (nn_759, nn_756, n_668);
  nand eco113 (nn_758, nn_143, nn_552);
  nand eco114 (nn_636, nn_634, nn_635);
  not eco115 (nwc35, n_472);
  not eco116 (nwc36, nn_547);
  nand eco117 (nn_547, nn_641, nn_642);
  not eco118 (nwc37, nn_369);
  nand eco119 (nn_369, n_490, nn_657);
  not eco120 (nwc38, nn_47);
  or eco121 (nn_652, nwc40, nn_524);
  not eco122 (nwc39, n_549);
  nand eco123 (nn_410, nn_521, nn_615);
  or eco124 (nn_642, nn_264, nn_410);
  or eco125 (nn_756, nwc42, nn_143);
  or eco126 (nn_634, nn_185, nn_56);
  or eco127 (nn_635, nn_264, nwc45);
  nand eco128 (nn_143, nn_521, n_474);
  or eco129 (nn_552, nn_597, nwc41);
  not eco130 (nwc40, nn_651);
  nand eco131 (nn_524, nn_455, n_534);
  nand eco132 (nn_651, nn_555, n_489);
  nand eco133 (nn_657, n_489, nn_410);
  nand eco134 (nn_662, nn_540, nn_56);
  nand eco135 (nn_597, nn_595, nn_596);
  not eco136 (nwc41, n_472);
  not eco137 (nwc42, nn_553);
  nand eco138 (nn_553, nn_602, nn_603);
  nand eco139 (nn_56, nn_620, n_665);
  nand eco140 (nn_611, nn_543, n_471);
  not eco141 (nwc43, nn_746);
  nand eco142 (nn_747, nn_744, n_683);
  nand eco143 (nn_746, n_573, nn_548);
  nand eco144 (nn_538, n_549, nn_627);
  or eco145 (nn_627, nn_626, nwc46);
  not eco146 (nwc44, nn_56);
  nand eco147 (nn_555, nn_521, nn_606);
  not eco148 (nwc45, nn_410);
  nand eco149 (nn_620, nn_539, nn_41);
  or eco150 (nn_602, nn_185, nwc49);
  or eco151 (nn_603, nn_264, nn_360);
  or eco152 (nn_744, nwc50, n_573);
  nand eco153 (nn_626, nn_537, n_535);
  not eco154 (nwc46, n_544);
  or eco155 (nn_595, nn_185, nn_41);
  or eco156 (nn_596, nn_264, nwc48);
  or eco157 (nn_521, wc1, \b[2]);
  nand eco158 (nn_615, n_474, nn_360);
  nand eco159 (nn_606, nn_554, n_474);
  or eco160 (nn_548, nn_570, nwc47);
  nand eco161 (nn_570, nn_568, nn_569);
  not eco162 (nwc47, n_472);
  nand eco163 (nn_41, nn_584, n_680);
  or eco164 (nn_612, n_471, n_582);
  or eco165 (nn_537, nn_524, nwc51);
  not eco166 (nwc48, nn_360);
  nand eco167 (nn_360, n_506, nn_579);
  not eco168 (nwc49, nn_41);
  not eco169 (nwc50, nn_549);
  nand eco170 (nn_549, nn_575, nn_576);
  nand eco171 (nn_554, n_506, nn_735);
  nand eco172 (nn_543, nn_496, nn_561);
  nand eco173 (nn_579, n_505, nn_496);
  not eco174 (nwc51, nn_588);
  nand eco175 (nn_588, n_482, nn_475);
  or eco176 (nn_735, nn_561, nwc55);
  or eco177 (nn_584, nwc52, n_582);
  or eco178 (nn_575, nn_185, n_582);
  or eco179 (nn_576, nn_264, nn_496);
  or eco180 (nn_568, nn_185, nwc53);
  or eco181 (nn_569, nn_264, nwc54);
  or eco182 (nn_561, wc47, \b[0]);
  not eco183 (nwc52, nn_541);
  not eco184 (nwc53, n_582);
  not eco185 (nwc54, nn_496);
  not eco186 (nwc55, n_505);
  not eco187 (nwc63, nn_69);
  not eco188 (nwc64, nn_711);
  not eco189 (nwc65, nn_69);
  not eco190 (nwc66, nn_69);
  not eco191 (nwc67, nn_69);
  not eco192 (nwc68, nn_69);
  not eco193 (nwc69, nn_69);
endmodule
// cost:187