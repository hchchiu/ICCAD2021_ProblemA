module top_eco(Gate);
  output Gate;
  assign Gate = 1'b0;
endmodule
