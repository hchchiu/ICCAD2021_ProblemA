module top(clk, oe, a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], b[0], b[1], b[2], b[3], b[4], b[5], b[6], b[7], op[0], op[1], y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7], parity, overflow, greater, is_eq, less);
  input clk, oe, a[0], a[1], a[2], a[3];
  input a[4], a[5], a[6], a[7], b[0], b[1];
  input b[2], b[3], b[4], b[5], b[6], b[7];
  input op[0], op[1];
  output y[0], y[1], y[2], y[3], y[4], y[5];
  output y[6], y[7], parity, overflow, greater, is_eq;
  output less;
  or eco1 (patchNew_n_368, patchNew_wc46, op[0]);
  not eco2 (patchNew_wc39, patchNew_n_121);
  nand eco3 (patchNew_n_249, patchNew_n_543, patchNew_n_544);
  or eco4 (patchNew_n_537, patchNew_wc31, n_551);
  or eco5 (patchNew_n_540, patchNew_sub_33_29_n_32, patchNew_sub_33_29_n_60);
  or eco6 (patchNew_n_536, patchNew_sub_33_29_n_48, n_551);
  nand eco7 (patchNew_n_535, patchNew_sub_33_29_n_48, n_551);
  nand eco8 (patchNew_n_382, patchNew_n_297, patchNew_n_121);
  nand eco9 (patchNew_n_499, patchNew_n_295, patchNew_sub_33_29_n_32);
  not eco10 (patchNew_gt_43_12_n_34, a[1]);
  or eco11 (patchNew_n_297, patchNew_n_364, patchNew_n_113);
  nand eco12 (parity, n_854, n_855);
  assign overflow = y[7];
  and eco14 (y[0], patchNew_temp_y0, patchNew_wc53);
  not eco15 (greater, patchNew_gt_43_12_n_36);
  and eco16 (y[1], patchNew_temp_y1, patchNew_wc52);
  and eco17 (y[2], patchNew_wc54, patchNew_temp_y2);
  and eco18 (y[3], patchNew_wc55, patchNew_temp_y3);
  and eco19 (y[4], patchNew_wc56, patchNew_temp_y4);
  and eco20 (y[5], patchNew_wc57, patchNew_temp_y5);
  nor eco21 (y[6], patchNew_n_472, patchNew_n_358);
  not eco22 (y[7], patchNew_n_358);
  and eco23 (is_eq, patchNew_gt_43_12_n_36, patchNew_lt_44_17_n_36);
  and eco24 (less, patchNew_gt_43_12_n_36, patchNew_wc51);
  or eco25 (n_523, wc, a[3]);
  not eco26 (wc, b[3]);
  or eco27 (n_568, wc1, a[7]);
  not eco28 (wc1, b[7]);
  or eco29 (n_522, wc3, a[4]);
  or eco30 (n_525, wc4, a[2]);
  not eco31 (wc3, b[4]);
  not eco32 (wc4, b[2]);
  or eco33 (n_534, wc6, a[5]);
  or eco34 (n_569, b[7], wc7);
  not eco35 (wc6, b[5]);
  or eco36 (n_570, wc8, a[6]);
  not eco37 (wc7, a[7]);
  or eco38 (n_571, b[6], wc9);
  not eco39 (wc8, b[6]);
  or eco40 (n_590, a[4], b[4]);
  not eco41 (wc9, a[6]);
  or eco42 (n_594, a[3], b[3]);
  or eco43 (n_854, patchNew_wc3, patchNew_n_110);
  or eco44 (n_596, a[2], b[2]);
  or eco45 (n_855, patchNew_n_241, patchNew_wc4);
  nand eco46 (n_558, n_534, n_535);
  or eco47 (n_535, wc58, b[5]);
  nand eco48 (n_545, n_521, n_522);
  or eco49 (n_531, wc56, b[3]);
  nand eco50 (n_554, n_523, n_531);
  or eco51 (n_521, wc57, b[4]);
  nand eco52 (n_739, a[4], b[4]);
  nand eco53 (n_718, a[3], b[3]);
  nand eco54 (n_577, n_535, n_571);
  nand eco55 (n_551, n_524, n_525);
  nand eco56 (n_593, n_569, n_682);
  or eco57 (n_682, n_681, wc42);
  or eco58 (n_524, wc55, b[2]);
  nand eco59 (n_676, a[2], b[2]);
  nand eco60 (n_681, n_592, n_568);
  not eco61 (wc42, n_570);
  or eco62 (n_592, n_577, wc47);
  nand eco63 (n_643, n_522, n_534);
  not eco64 (wc47, n_643);
  or eco65 (n_539, wc53, op[0]);
  nand eco66 (n_780, a[5], b[5]);
  not eco67 (wc53, op[1]);
  not eco68 (wc52, a[0]);
  not eco69 (wc54, a[1]);
  not eco70 (wc55, a[2]);
  not eco71 (wc57, a[4]);
  not eco72 (wc56, a[3]);
  not eco73 (wc58, a[5]);
  not eco74 (patchNew_wc31, patchNew_add_28_29_n_41);
  or eco75 (patchNew_n_541, patchNew_wc34, patchNew_add_28_29_n_53);
  or eco76 (patchNew_n_542, patchNew_add_28_29_n_21, patchNew_wc35);
  not eco77 (patchNew_wc34, patchNew_add_28_29_n_21);
  nand eco78 (patchNew_add_28_29_n_53, patchNew_n_296, patchNew_n_325);
  not eco79 (patchNew_wc35, patchNew_add_28_29_n_53);
  or eco80 (patchNew_n_538, patchNew_add_28_29_n_41, patchNew_wc32);
  nand eco81 (patchNew_n_381, patchNew_n_298, patchNew_gt_43_12_n_34);
  nand eco82 (patchNew_n_259, patchNew_n_541, patchNew_n_542);
  nand eco83 (patchNew_n_394, patchNew_sub_33_29_n_48, n_525);
  nand eco84 (patchNew_n_539, patchNew_sub_33_29_n_32, patchNew_sub_33_29_n_60);
  nand eco85 (patchNew_n_397, patchNew_add_28_29_n_41, n_596);
  or eco86 (patchNew_n_276, b[5], wc58);
  or eco87 (patchNew_n_502, patchNew_wc36, patchNew_add_28_29_n_21);
  nand eco88 (patchNew_n_243, patchNew_n_537, patchNew_n_538);
  or eco89 (patchNew_lt_44_17_n_44, wc55, b[2]);
  nand eco90 (patchNew_n_375, patchNew_n_292, a[1]);
  or eco91 (patchNew_n_376, patchNew_wc37, patchNew_n_121);
  nand eco92 (patchNew_sub_33_29_n_32, patchNew_lt_44_17_n_37, patchNew_n_113);
  or eco93 (patchNew_n_318, patchNew_n_121, wc54);
  not eco94 (patchNew_wc37, patchNew_n_359);
  not eco95 (patchNew_wc36, patchNew_n_296);
  nand eco96 (patchNew_sub_33_29_n_60, patchNew_n_318, patchNew_n_295);
  nand eco97 (patchNew_n_325, patchNew_n_121, a[1]);
  not eco98 (patchNew_wc32, n_551);
  not eco99 (patchNew_wc46, a[1]);
  or eco100 (patchNew_n_543, patchNew_wc40, patchNew_n_121);
  or eco101 (patchNew_n_544, a[1], patchNew_wc41);
  nand eco102 (patchNew_n_364, a[1], a[0]);
  or eco103 (patchNew_n_330, n_539, patchNew_wc44);
  or eco104 (patchNew_n_331, patchNew_wc43, a[0]);
  or eco105 (patchNew_n_359, patchNew_n_363, patchNew_wc42);
  or eco106 (patchNew_n_363, a[1], a[0]);
  not eco107 (patchNew_wc42, patchNew_n_113);
  not eco108 (patchNew_wc40, a[1]);
  not eco109 (patchNew_wc41, patchNew_n_121);
  nand eco110 (patchNew_n_320, n_739, n_780);
  or eco111 (patchNew_n_317, n_521, patchNew_wc58);
  not eco112 (patchNew_wc58, n_534);
  nand eco113 (patchNew_gt_43_12_n_36, n_593, patchNew_n_445);
  or eco114 (patchNew_n_472, patchNew_wc17, op[1]);
  or eco115 (patchNew_n_358, patchNew_n_468, patchNew_n_469);
  not eco116 (patchNew_wc51, patchNew_lt_44_17_n_36);
  nand eco117 (patchNew_temp_y0, patchNew_n_390, patchNew_n_391);
  not eco118 (patchNew_wc53, patchNew_n_358);
  nand eco119 (patchNew_temp_y1, patchNew_n_438, patchNew_n_439);
  not eco120 (patchNew_wc52, patchNew_n_358);
  not eco121 (patchNew_wc54, patchNew_n_358);
  nand eco122 (patchNew_temp_y2, patchNew_n_462, patchNew_n_463);
  not eco123 (patchNew_wc55, patchNew_n_358);
  nand eco124 (patchNew_temp_y3, patchNew_n_483, patchNew_n_484);
  not eco125 (patchNew_wc56, patchNew_n_358);
  nand eco126 (patchNew_temp_y4, patchNew_n_489, patchNew_n_490);
  not eco127 (patchNew_wc57, patchNew_n_358);
  nand eco128 (patchNew_temp_y5, patchNew_n_495, patchNew_n_496);
  nand eco129 (patchNew_lt_44_17_n_36, patchNew_lt_44_17_n_88, patchNew_n_442);
  not eco130 (patchNew_wc3, patchNew_n_241);
  nand eco131 (patchNew_n_110, patchNew_n_508, patchNew_n_509);
  nand eco132 (patchNew_n_241, patchNew_n_505, patchNew_n_506);
  not eco133 (patchNew_wc4, patchNew_n_110);
  or eco134 (patchNew_n_390, patchNew_n_389, patchNew_n_113);
  nand eco135 (patchNew_n_391, patchNew_n_280, patchNew_n_113);
  or eco136 (patchNew_n_438, op[1], patchNew_wc25);
  nand eco137 (patchNew_n_439, patchNew_n_290, op[1]);
  or eco138 (patchNew_n_462, op[1], patchNew_wc23);
  nand eco139 (patchNew_n_463, patchNew_n_286, op[1]);
  or eco140 (patchNew_n_483, op[1], patchNew_wc15);
  nand eco141 (patchNew_n_484, patchNew_n_282, op[1]);
  or eco142 (patchNew_n_489, op[1], patchNew_wc14);
  nand eco143 (patchNew_n_490, patchNew_n_288, op[1]);
  or eco144 (patchNew_n_495, op[1], patchNew_wc13);
  nand eco145 (patchNew_n_496, patchNew_n_284, op[1]);
  nand eco146 (patchNew_n_445, patchNew_n_300, patchNew_gt_43_12_n_87);
  nand eco147 (patchNew_lt_44_17_n_88, patchNew_n_346, patchNew_n_347);
  nand eco148 (patchNew_n_442, patchNew_n_294, patchNew_lt_44_17_n_87);
  or eco149 (patchNew_n_508, patchNew_wc7, patchNew_n_109);
  or eco150 (patchNew_n_509, patchNew_n_242, patchNew_wc8);
  or eco151 (patchNew_n_505, patchNew_wc5, patchNew_temp_y5);
  or eco152 (patchNew_n_506, patchNew_temp_y0, patchNew_wc6);
  nand eco153 (patchNew_add_28_29_n_21, a[0], patchNew_n_113);
  nand eco154 (patchNew_n_113, patchNew_n_306, patchNew_n_360);
  or eco155 (patchNew_n_306, wc8, clk);
  nand eco156 (patchNew_n_360, b[0], clk);
  not eco157 (patchNew_wc17, patchNew_n_278);
  or eco158 (patchNew_n_468, patchNew_wc65, op[1]);
  nand eco159 (patchNew_n_469, op[0], patchNew_lt_44_17_n_68);
  not eco160 (patchNew_wc7, patchNew_n_242);
  nand eco161 (patchNew_n_242, patchNew_n_510, patchNew_n_511);
  or eco162 (patchNew_n_510, patchNew_wc9, patchNew_temp_y1);
  or eco163 (patchNew_n_511, patchNew_temp_y4, patchNew_wc10);
  nand eco164 (patchNew_n_292, patchNew_n_113, patchNew_lt_44_17_n_37);
  not eco165 (patchNew_lt_44_17_n_37, a[0]);
  or eco166 (patchNew_n_295, patchNew_wc0, a[1]);
  not eco167 (patchNew_wc0, patchNew_n_121);
  nand eco168 (patchNew_n_121, patchNew_n_361, patchNew_n_362);
  or eco169 (patchNew_n_296, patchNew_n_121, a[1]);
  or eco170 (patchNew_n_361, wc1, clk);
  nand eco171 (patchNew_n_362, b[1], clk);
  or eco172 (patchNew_n_298, patchNew_n_113, wc52);
  nand eco173 (patchNew_n_301, patchNew_sub_33_29_n_54, patchNew_lt_44_17_n_71);
  nand eco174 (patchNew_sub_33_29_n_54, patchNew_lt_44_17_n_66, patchNew_n_412);
  not eco175 (patchNew_lt_44_17_n_71, patchNew_n_262);
  nand eco176 (patchNew_lt_44_17_n_66, patchNew_n_24, n_523);
  nand eco177 (patchNew_n_412, patchNew_sub_33_29_n_48, patchNew_lt_44_17_n_65);
  nand eco178 (patchNew_n_262, n_522, n_534);
  nand eco179 (patchNew_n_24, n_531, patchNew_lt_44_17_n_44);
  nand eco180 (patchNew_sub_33_29_n_48, patchNew_n_318, patchNew_n_499);
  not eco181 (patchNew_lt_44_17_n_65, patchNew_n_27);
  not eco182 (patchNew_wc5, patchNew_temp_y0);
  not eco183 (patchNew_wc6, patchNew_temp_y5);
  nand eco184 (patchNew_n_109, patchNew_n_513, patchNew_n_514);
  not eco185 (patchNew_wc8, patchNew_n_109);
  not eco186 (patchNew_wc9, patchNew_temp_y4);
  not eco187 (patchNew_wc13, patchNew_n_283);
  nand eco188 (patchNew_n_284, patchNew_n_342, patchNew_n_343);
  nand eco189 (patchNew_n_389, a[0], n_539);
  nand eco190 (patchNew_n_280, patchNew_n_330, patchNew_n_331);
  nand eco191 (patchNew_n_283, patchNew_n_477, patchNew_n_478);
  or eco192 (patchNew_n_342, op[0], n_780);
  nand eco193 (patchNew_n_343, n_558, op[0]);
  or eco194 (patchNew_n_513, patchNew_wc11, patchNew_temp_y2);
  or eco195 (patchNew_n_514, patchNew_temp_y3, patchNew_wc12);
  nand eco196 (patchNew_n_426, patchNew_add_28_29_n_47, patchNew_add_28_29_n_50);
  nand eco197 (patchNew_add_28_29_n_47, patchNew_add_28_29_n_45, patchNew_n_415);
  and eco198 (patchNew_add_28_29_n_50, patchNew_n_312, n_590);
  nand eco199 (patchNew_add_28_29_n_45, n_594, patchNew_n_323);
  nand eco200 (patchNew_n_415, patchNew_add_28_29_n_41, patchNew_add_28_29_n_44);
  or eco201 (patchNew_n_312, b[5], a[5]);
  nand eco202 (patchNew_n_258, patchNew_n_533, patchNew_n_534);
  nand eco203 (patchNew_n_533, patchNew_sub_33_29_n_63, n_554);
  or eco204 (patchNew_n_534, patchNew_sub_33_29_n_63, n_554);
  nand eco205 (patchNew_sub_33_29_n_63, patchNew_lt_44_17_n_44, patchNew_n_394);
  not eco206 (patchNew_wc25, patchNew_n_289);
  nand eco207 (patchNew_n_289, patchNew_n_402, patchNew_n_403);
  not eco208 (patchNew_wc11, patchNew_temp_y3);
  not eco209 (patchNew_wc12, patchNew_temp_y2);
  not eco210 (patchNew_wc10, patchNew_temp_y1);
  nand eco211 (patchNew_n_290, patchNew_n_369, patchNew_n_370);
  not eco212 (patchNew_wc14, patchNew_n_287);
  nand eco213 (patchNew_n_288, patchNew_n_354, patchNew_n_355);
  or eco214 (patchNew_n_477, patchNew_wc16, op[0]);
  nand eco215 (patchNew_n_478, patchNew_n_253, op[0]);
  not eco216 (patchNew_wc16, patchNew_n_252);
  nand eco217 (patchNew_n_253, patchNew_n_521, patchNew_n_522);
  not eco218 (patchNew_wc23, patchNew_n_285);
  nand eco219 (patchNew_n_286, patchNew_n_348, patchNew_n_349);
  not eco220 (patchNew_wc15, patchNew_n_281);
  nand eco221 (patchNew_n_282, patchNew_n_336, patchNew_n_337);
  nand eco222 (patchNew_n_287, patchNew_n_456, patchNew_n_457);
  nand eco223 (patchNew_n_281, patchNew_n_450, patchNew_n_451);
  or eco224 (patchNew_n_336, op[0], n_718);
  nand eco225 (patchNew_n_337, n_554, op[0]);
  or eco226 (patchNew_n_456, patchNew_wc20, op[0]);
  nand eco227 (patchNew_n_457, patchNew_n_255, op[0]);
  not eco228 (patchNew_wc20, patchNew_n_254);
  nand eco229 (patchNew_n_255, patchNew_n_531, patchNew_n_532);
  or eco230 (patchNew_n_354, op[0], n_739);
  nand eco231 (patchNew_n_355, n_545, op[0]);
  nand eco232 (patchNew_n_252, patchNew_n_524, patchNew_n_525);
  nand eco233 (patchNew_n_521, patchNew_sub_33_29_n_67, n_558);
  or eco234 (patchNew_n_522, patchNew_sub_33_29_n_67, n_558);
  nand eco235 (patchNew_sub_33_29_n_67, n_521, patchNew_n_418);
  or eco236 (patchNew_n_524, patchNew_wc18, n_558);
  or eco237 (patchNew_n_525, patchNew_add_28_29_n_60, patchNew_wc19);
  or eco238 (patchNew_n_450, patchNew_wc21, op[0]);
  nand eco239 (patchNew_n_451, patchNew_n_258, op[0]);
  not eco240 (patchNew_wc21, patchNew_n_257);
  nand eco241 (patchNew_n_254, patchNew_n_529, patchNew_n_530);
  not eco242 (patchNew_wc18, patchNew_add_28_29_n_60);
  nand eco243 (patchNew_add_28_29_n_60, n_739, patchNew_n_421);
  not eco244 (patchNew_wc19, n_558);
  or eco245 (patchNew_n_278, patchNew_wc22, patchNew_n_427);
  not eco246 (patchNew_wc22, patchNew_n_426);
  or eco247 (patchNew_n_427, patchNew_wc45, op[0]);
  not eco248 (patchNew_wc45, patchNew_add_28_29_n_51);
  nand eco249 (patchNew_n_531, patchNew_sub_33_29_n_54, n_545);
  or eco250 (patchNew_n_532, patchNew_sub_33_29_n_54, n_545);
  nand eco251 (patchNew_n_257, patchNew_n_527, patchNew_n_528);
  nand eco252 (patchNew_n_418, patchNew_sub_33_29_n_54, n_522);
  nand eco253 (patchNew_n_421, patchNew_add_28_29_n_47, n_590);
  or eco254 (patchNew_n_529, patchNew_wc28, n_545);
  or eco255 (patchNew_n_530, patchNew_add_28_29_n_47, patchNew_wc66);
  nand eco256 (patchNew_n_285, patchNew_n_432, patchNew_n_433);
  or eco257 (patchNew_n_348, op[0], n_676);
  nand eco258 (patchNew_n_349, n_551, op[0]);
  not eco259 (patchNew_wc65, patchNew_n_301);
  not eco260 (patchNew_lt_44_17_n_68, patchNew_n_34);
  nand eco261 (patchNew_n_34, patchNew_n_317, patchNew_n_276);
  or eco262 (patchNew_n_527, patchNew_wc26, n_554);
  or eco263 (patchNew_n_528, patchNew_add_28_29_n_56, patchNew_wc27);
  not eco264 (patchNew_wc28, patchNew_add_28_29_n_47);
  not eco265 (patchNew_wc66, n_545);
  not eco266 (patchNew_wc26, patchNew_add_28_29_n_56);
  nand eco267 (patchNew_add_28_29_n_56, n_676, patchNew_n_397);
  not eco268 (patchNew_wc27, n_554);
  or eco269 (patchNew_n_346, patchNew_n_34, patchNew_n_308);
  nand eco270 (patchNew_n_347, n_569, patchNew_n_307);
  nand eco271 (patchNew_n_294, patchNew_lt_44_17_n_66, patchNew_n_406);
  nor eco272 (patchNew_lt_44_17_n_87, patchNew_n_262, patchNew_n_307);
  nand eco273 (patchNew_n_300, patchNew_gt_43_12_n_66, patchNew_n_409);
  nor eco274 (patchNew_gt_43_12_n_87, patchNew_n_332, patchNew_n_308);
  nand eco275 (patchNew_n_308, n_569, n_571);
  nand eco276 (patchNew_n_307, n_568, n_570);
  nand eco277 (patchNew_n_406, patchNew_n_293, patchNew_lt_44_17_n_65);
  nand eco278 (patchNew_add_28_29_n_51, patchNew_n_312, patchNew_n_320);
  not eco279 (patchNew_wc44, a[0]);
  not eco280 (patchNew_wc43, n_539);
  or eco281 (patchNew_n_369, patchNew_n_368, patchNew_wc39);
  nand eco282 (patchNew_n_370, patchNew_n_249, op[0]);
  or eco283 (patchNew_n_432, patchNew_wc67, op[0]);
  nand eco284 (patchNew_n_433, patchNew_n_244, op[0]);
  not eco285 (patchNew_wc67, patchNew_n_243);
  nand eco286 (patchNew_n_244, patchNew_n_535, patchNew_n_536);
  nand eco287 (patchNew_gt_43_12_n_66, patchNew_n_27, n_531);
  nand eco288 (patchNew_n_409, patchNew_n_299, patchNew_gt_43_12_n_65);
  nand eco289 (patchNew_n_332, n_521, patchNew_n_276);
  nand eco290 (patchNew_n_293, patchNew_n_375, patchNew_n_376);
  nand eco291 (patchNew_n_323, n_676, n_718);
  nand eco292 (patchNew_add_28_29_n_41, patchNew_n_325, patchNew_n_502);
  and eco293 (patchNew_add_28_29_n_44, n_594, n_596);
  or eco294 (patchNew_n_402, patchNew_wc30, op[0]);
  nand eco295 (patchNew_n_403, patchNew_n_260, op[0]);
  not eco296 (patchNew_wc30, patchNew_n_259);
  nand eco297 (patchNew_n_260, patchNew_n_539, patchNew_n_540);
  nand eco298 (patchNew_n_27, n_523, n_525);
  nand eco299 (patchNew_n_299, patchNew_n_381, patchNew_n_382);
  not eco300 (patchNew_gt_43_12_n_65, patchNew_n_24);
endmodule