module top_eco(g4671, g4672, g4669, g4705, g4706, g4707, g4708, g4674, g4676, g4677, g4680, g4681, g4682, g4683, g4684, g4685, g4687, g4688, g4689, g4691, g4692, g4693, g4694, g4695, g4696, g4697, g4698, g4699, g4700, g4701, g4703, g4704, g471, g4709, g4710, g4711, g4715, g4716, g4717, g4718, g4719, g4720, g4721, g4725, g4726, g4727, g4729, g4731, g4732, g4735, g4736, g4738, g4740, g4741, g4743, g4744, g4746, g4748, g4749, g4750, g4751, g4752, g4753, g4754, g4755, g4756, g4757, g4758, g4764, g4766, g4767, g4768, g4769, g4770, g4771, g4772, g4773, g4774, g4775, g4776, g4778, g4779, g4780, g4781, g4782, g4784, g4785, g4787, g4788, g4789, g4790, g4791, g4793, g4794, g4795, g4796, g4797, g4798, g4799, g4800, g4802, g4803, g4806, g4807, g4808, g4809, g4810, g4811, g4812, g4813, g4814, g4815, g1357, g1240, g923, g445, g448, g450, g454, g460, g461, g476, g478, g483, g487, g491, g492, g495, g497, g501, g505, g509, g510, g511_g4785_96, g518, g533, g535, g536, g538, g542, g550, g553, g555, g569, g575, g576, g580, g581, g582, g593, g600, g608, g609, g610, g618, g624, g625, g627, g630, g632, g633, g643, g648, g658, g665, g670, g685, g686, g687, g688, g703, g705, g706, g710, g720, g724, g730, g731, g739, g750, g753, g760, g771, g790, g801, g804, g813, g839, g864, g878, g904, g953, g987, g1015, g1024, g1035, g1049, g4702_g4785_189, g1062, g1068, g1122, g1123, g1156, g1171, g1308, g1332, g1340, g4849, g4851, g4852, g4853, g4854, g4855, g4856, g4857, g4861, g4862, g4863, g4864, g4865, g4866, g4867, g4868, g4869, g4870, g4871, g4873, g4874, g4879, g4880, g4881, g4882, g4883, g4884, g4886, g4888, g4889, g992, g1350, g1358, g991, g983, g1352, g989, g1343, g1325, g1339);
  input g4671, g4672, g4669, g4705;
  input g4706, g4707, g4708, g4674, g4676;
  input g4677, g4680, g4681, g4682, g4683;
  input g4684, g4685, g4687, g4688, g4689;
  input g4691, g4692, g4693, g4694, g4695;
  input g4696, g4697, g4698, g4699, g4700;
  input g4701, g4703, g4704, g471, g4709;
  input g4710, g4711, g4715, g4716, g4717;
  input g4718, g4719, g4720, g4721, g4725;
  input g4726, g4727, g4729, g4731, g4732;
  input g4735, g4736, g4738, g4740, g4741;
  input g4743, g4744, g4746, g4748, g4749;
  input g4750, g4751, g4752, g4753, g4754;
  input g4755, g4756, g4757, g4758, g4764;
  input g4766, g4767, g4768, g4769, g4770;
  input g4771, g4772, g4773, g4774, g4775;
  input g4776, g4778, g4779, g4780, g4781;
  input g4782, g4784, g4785, g4787, g4788;
  input g4789, g4790, g4791, g4793, g4794;
  input g4795, g4796, g4797, g4798, g4799;
  input g4800, g4802, g4803, g4806, g4807;
  input g4808, g4809, g4810, g4811, g4812;
  input g4813, g4814, g4815, g1357, g1240;
  input g923, g445, g448, g450, g454;
  input g460, g461, g476, g478, g483;
  input g487, g491, g492, g495, g497;
  input g501, g505, g509, g510, g511_g4785_96;
  input g518, g533, g535, g536, g538;
  input g542, g550, g553, g555, g569;
  input g575, g576, g580, g581, g582;
  input g593, g600, g608, g609, g610;
  input g618, g624, g625, g627, g630;
  input g632, g633, g643, g648, g658;
  input g665, g670, g685, g686, g687;
  input g688, g703, g705, g706, g710;
  input g720, g724, g730, g731, g739;
  input g750, g753, g760, g771, g790;
  input g801, g804, g813, g839, g864;
  input g878, g904, g953, g987, g1015;
  input g1024, g1035, g1049, g4702_g4785_189, g1062;
  input g1068, g1122, g1123, g1156, g1171;
  input g1308, g1332, g1340;
  output g4849, g4851, g4852, g4853;
  output g4854, g4855, g4856, g4857, g4861;
  output g4862, g4863, g4864, g4865, g4866;
  output g4867, g4868, g4869, g4870, g4871;
  output g4873, g4874, g4879, g4880, g4881;
  output g4882, g4883, g4884, g4886, g4888;
  output g4889, g992, g1350, g1358, g991;
  output g983, g1352, g989, g1343, g1325;
  output g1339;
  buf eco1 (g4849, patchNew_n1040);
  buf eco2 (g4851, patchNew_n593);
  buf eco3 (g4852, patchNew_n477);
  buf eco4 (g4853, patchNew_n1037);
  buf eco5 (g4854, patchNew_n747);
  buf eco6 (g4855, patchNew_n770);
  buf eco7 (g4856, patchNew_n1031);
  buf eco8 (g4857, patchNew_n373);
  buf eco9 (g4861, patchNew_n244);
  buf eco10 (g4862, patchNew_n378);
  buf eco11 (g4863, patchNew_n1034);
  buf eco12 (g4864, patchNew_n400);
  buf eco13 (g4865, patchNew_n348);
  buf eco14 (g4866, patchNew_n448);
  buf eco15 (g4867, patchNew_n494);
  buf eco16 (g4868, patchNew_n1029);
  buf eco17 (g4869, patchNew_n1029);
  buf eco18 (g4870, patchNew_n1033);
  buf eco19 (g4871, patchNew_n1033);
  buf eco20 (g4873, patchNew_n1026);
  buf eco21 (g4874, patchNew_n1026);
  buf eco22 (g4879, patchNew_n976);
  buf eco23 (g4880, patchNew_n977);
  buf eco24 (g4881, patchNew_n1017);
  buf eco25 (g4882, patchNew_n1001);
  buf eco26 (g4883, patchNew_n1000);
  buf eco27 (g4884, patchNew_n1000);
  buf eco28 (g4886, patchNew_n588);
  buf eco29 (g4888, patchNew_n837);
  buf eco30 (g4889, patchNew_n838);
  nand eco31 (g992, patchNew_n139_n140_84_n141_85, g4810);
  nand eco32 (g1350, patchNew_n1043, g4787);
  nand eco33 (g1358, patchNew_n1045, g4815);
  not eco34 (g991, patchNew_n1040);
  nand eco35 (g983, g4790, patchNew_n321);
  nand eco36 (g1352, patchNew_n116_n121_79_n28_80, patchNew_n593);
  nand eco37 (g989, patchNew_n121_n1038_81_n116_82, patchNew_n593);
  nand eco38 (g1343, patchNew_n1021, patchNew_n1022);
  nand eco39 (g1325, patchNew_1'b1_n1018_78, patchNew__xnor_GATE_0);
  not eco40 (g1339, patchNew_n835);
  and eco41 (patchNew_n1040, patchNew_new_n263_, patchNew_new_n266_);
  nor eco42 (patchNew_n593, patchNew_new_n268_, patchNew_new_n269_);
  and eco43 (patchNew_n477, patchNew__not_GATE_9, patchNew_new_n277_);
  nor eco44 (patchNew_n1037, patchNew_new_n282_, patchNew_new_n286_);
  nor eco45 (patchNew_n747, patchNew_new_n289_, patchNew_new_n296_);
  and eco46 (patchNew_n770, patchNew__not_GATE_17, patchNew_new_n305_);
  nor eco47 (patchNew_n1031, patchNew_new_n313_, patchNew_new_n314_);
  and eco48 (patchNew_n373, patchNew__not_GATE_23, patchNew_new_n324_);
  or eco49 (patchNew_n244, patchNew_new_n328_, patchNew__not_GATE_27);
  or eco50 (patchNew_n378, patchNew_new_n323_, patchNew_new_n333_);
  not eco51 (patchNew_n1034, patchNew_n1031);
  not eco52 (patchNew_n400, patchNew_n770);
  or eco53 (patchNew_n348, patchNew_new_n339_, patchNew_new_n341_);
  or eco54 (patchNew_n448, patchNew_new_n344_, patchNew__not_GATE_32);
  or eco55 (patchNew_n494, patchNew__not_GATE_33, patchNew_new_n352_);
  or eco56 (patchNew_n1029, patchNew_new_n365_, patchNew_new_n366_);
  or eco57 (patchNew_n1033, patchNew_new_n368_, patchNew_new_n369_);
  or eco58 (patchNew_n1026, patchNew_new_n372_, patchNew_new_n382_);
  and eco59 (patchNew_n976, patchNew__not_GATE_86, patchNew_new_n532_);
  not eco60 (patchNew_n977, patchNew_n976);
  nor eco61 (patchNew_n1017, patchNew_new_n548_, patchNew_new_n551_);
  and eco62 (patchNew_n1001, patchNew__not_GATE_110, patchNew_new_n583_);
  or eco63 (patchNew_n1000, patchNew_new_n585_, patchNew_new_n609_);
  or eco64 (patchNew_n588, patchNew_new_n638_, patchNew_new_n701_);
  and eco65 (patchNew_n837, patchNew__not_GATE_179, patchNew_new_n721_);
  not eco66 (patchNew_n838, patchNew_n837);
  and eco67 (patchNew_n321, patchNew__not_GATE_41, patchNew_new_n380_);
  nor eco68 (patchNew_new_n308_, g4785, patchNew_new_n307_);
  and eco69 (patchNew_new_n320_, g670, patchNew__not_GATE_21);
  or eco70 (patchNew_n835, patchNew_new_n715_, patchNew__not_GATE_177);
  buf eco71 (patchNew_1'b1_n1018_78, g4812);
  or eco72 (patchNew_n1021, g4790, patchNew_new_n371_);
  or eco73 (patchNew_n1022, g864, patchNew_new_n364_);
  nand eco74 (patchNew_n116_n121_79_n28_80, g987, g4696);
  or eco75 (patchNew_n121_n1038_81_n116_82, patchNew__not_GATE_183, patchNew_new_n730_);
  not eco76 (patchNew_n1043, g1357);
  buf eco77 (patchNew_n1045, patchNew_n1043);
  or eco78 (patchNew_n139_n140_84_n141_85, patchNew__not_GATE_184, patchNew_new_n732_);
  not eco79 (patchNew_n1050, g706);
  xnor eco80 (patchNew__xnor_GATE_3, patchNew_new_n574_, patchNew_new_n511_);
  xnor eco81 (patchNew__xnor_GATE_4, patchNew_new_n587_, patchNew_new_n593_);
  xnor eco82 (patchNew__xnor_GATE_5, patchNew_n348, patchNew_n494);
  xnor eco83 (patchNew__xnor_GATE_6, g4809, patchNew_new_n486_);
  xnor eco84 (patchNew__xnor_GATE_7, g4793, patchNew_new_n493_);
  xnor eco85 (patchNew__xnor_GATE_8, patchNew_n477, patchNew_n1037);
  xnor eco86 (patchNew__xnor_GATE_9, patchNew_new_n371_, patchNew_new_n535_);
  xnor eco87 (patchNew__xnor_GATE_10, patchNew_n770, patchNew_new_n659_);
  xnor eco88 (patchNew__xnor_GATE_11, patchNew_new_n705_, patchNew_new_n710_);
  and eco89 (patchNew_new_n562_, g1122, g4752);
  and eco90 (patchNew_new_n563_, g4782, g501);
  and eco91 (patchNew_new_n564_, g4772, g706);
  and eco92 (patchNew_new_n565_, patchNew__not_GATE_102, g497);
  not eco93 (patchNew__not_GATE_102, g1156);
  nor eco94 (patchNew_new_n566_, patchNew_new_n563_, patchNew_new_n564_);
  and eco95 (patchNew_new_n567_, patchNew__not_GATE_103, patchNew_new_n566_);
  not eco96 (patchNew__not_GATE_103, patchNew_new_n565_);
  nor eco97 (patchNew_new_n568_, patchNew_new_n562_, patchNew_new_n567_);
  and eco98 (patchNew_new_n572_, patchNew_new_n568_, patchNew__xnor_GATE_2);
  nor eco99 (patchNew_new_n573_, patchNew_new_n568_, patchNew__xnor_GATE_2);
  nor eco100 (patchNew_new_n574_, patchNew_new_n572_, patchNew_new_n573_);
  and eco101 (patchNew_new_n578_, patchNew__xnor_GATE_1, patchNew__xnor_GATE_3);
  nor eco102 (patchNew_new_n579_, patchNew__xnor_GATE_1, patchNew__xnor_GATE_3);
  nor eco103 (patchNew_new_n580_, patchNew_new_n578_, patchNew_new_n579_);
  and eco104 (patchNew_new_n581_, patchNew__not_GATE_108, patchNew_new_n580_);
  not eco105 (patchNew__not_GATE_108, patchNew_new_n558_);
  and eco106 (patchNew_new_n582_, patchNew_new_n558_, patchNew__not_GATE_109);
  not eco107 (patchNew__not_GATE_109, patchNew_new_n580_);
  nor eco108 (patchNew_new_n583_, g4697, patchNew_new_n581_);
  not eco109 (patchNew__not_GATE_110, patchNew_new_n582_);
  nor eco110 (patchNew_new_n585_, g4791, patchNew_new_n547_);
  and eco111 (patchNew_new_n586_, patchNew__not_GATE_111, patchNew_new_n547_);
  not eco112 (patchNew__not_GATE_111, patchNew_new_n490_);
  nor eco113 (patchNew_new_n587_, patchNew_n321, patchNew_new_n586_);
  and eco114 (patchNew_new_n588_, patchNew_n244, patchNew_new_n371_);
  and eco115 (patchNew_new_n589_, patchNew_n244, patchNew_new_n364_);
  nor eco116 (patchNew_new_n590_, patchNew_n244, patchNew_new_n364_);
  nor eco117 (patchNew_new_n591_, patchNew_new_n589_, patchNew_new_n590_);
  and eco118 (patchNew_new_n592_, patchNew__not_GATE_112, patchNew_new_n591_);
  not eco119 (patchNew__not_GATE_112, patchNew_new_n371_);
  nor eco120 (patchNew_new_n593_, patchNew_new_n588_, patchNew_new_n592_);
  and eco121 (patchNew_new_n597_, patchNew_n770, patchNew_n448);
  nor eco122 (patchNew_new_n598_, patchNew_n770, patchNew_n448);
  nor eco123 (patchNew_new_n599_, patchNew_new_n597_, patchNew_new_n598_);
  and eco124 (patchNew_new_n603_, patchNew_new_n599_, patchNew__xnor_GATE_5);
  nor eco125 (patchNew_new_n604_, patchNew_new_n599_, patchNew__xnor_GATE_5);
  nor eco126 (patchNew_new_n605_, patchNew_new_n603_, patchNew_new_n604_);
  and eco127 (patchNew_new_n606_, patchNew__not_GATE_117, patchNew_new_n605_);
  not eco128 (patchNew__not_GATE_117, patchNew__xnor_GATE_4);
  and eco129 (patchNew_new_n607_, patchNew__not_GATE_118, patchNew__xnor_GATE_4);
  not eco130 (patchNew__not_GATE_118, patchNew_new_n605_);
  nor eco131 (patchNew_new_n608_, g1015, patchNew_new_n606_);
  and eco132 (patchNew_new_n609_, patchNew__not_GATE_119, patchNew_new_n608_);
  not eco133 (patchNew__not_GATE_119, patchNew_new_n607_);
  and eco134 (patchNew_new_n611_, patchNew__not_GATE_120, g760);
  not eco135 (patchNew__not_GATE_120, g1171);
  nor eco136 (patchNew_new_n612_, patchNew_new_n289_, patchNew_new_n611_);
  and eco137 (patchNew_new_n613_, patchNew__not_GATE_121, patchNew_new_n612_);
  not eco138 (patchNew__not_GATE_121, patchNew_new_n295_);
  and eco139 (patchNew_new_n614_, g4698, patchNew_n477);
  and eco140 (patchNew_new_n615_, g839, patchNew__not_GATE_122);
  not eco141 (patchNew__not_GATE_122, patchNew_new_n613_);
  and eco142 (patchNew_new_n616_, patchNew_new_n614_, patchNew_new_n615_);
  nor eco143 (patchNew_new_n617_, patchNew_new_n401_, patchNew_new_n616_);
  nor eco144 (patchNew_new_n618_, g4795, patchNew_new_n613_);
  and eco145 (patchNew_new_n301_, g4788, g4704);
  nor eco146 (patchNew_new_n300_, g801, g730);
  and eco147 (patchNew_new_n303_, patchNew_new_n301_, patchNew_new_n302_);
  and eco148 (patchNew_new_n279_, g4814, g4756);
  and eco149 (patchNew_new_n398_, g4773, g471);
  not eco150 (patchNew__not_GATE_10, patchNew_new_n281_);
  and eco151 (patchNew_new_n341_, g625, patchNew__not_GATE_30);
  and eco152 (patchNew_new_n497_, patchNew__not_GATE_72, patchNew_new_n496_);
  nor eco153 (patchNew_new_n517_, patchNew_new_n515_, patchNew_new_n516_);
  not eco154 (patchNew__not_GATE_72, patchNew_new_n470_);
  and eco155 (patchNew_new_n440_, g4672, g460);
  nor eco156 (patchNew_new_n441_, patchNew_new_n439_, patchNew_new_n440_);
  not eco157 (patchNew__not_GATE_27, patchNew_new_n330_);
  and eco158 (patchNew_new_n261_, g4721, g4754);
  not eco159 (patchNew__not_GATE_15, patchNew_new_n298_);
  and eco160 (patchNew_new_n302_, g878, g4725);
  and eco161 (patchNew_new_n326_, g4785, g4707);
  nor eco162 (patchNew_new_n333_, patchNew_new_n321_, patchNew_new_n332_);
  and eco163 (patchNew_new_n298_, g1024, g4736);
  not eco164 (patchNew__not_GATE_1, patchNew_new_n262_);
  and eco165 (patchNew_new_n299_, g625, patchNew__not_GATE_15);
  not eco166 (patchNew__not_GATE_39, patchNew_new_n374_);
  and eco167 (patchNew_new_n376_, g4788, g4699);
  not eco168 (patchNew__not_GATE_0, patchNew_new_n261_);
  and eco169 (patchNew_new_n276_, g610, g608);
  nor eco170 (patchNew_new_n324_, patchNew_new_n316_, patchNew_new_n323_);
  nor eco171 (patchNew_new_n365_, g4791, patchNew_new_n364_);
  nor eco172 (patchNew_new_n349_, g4785, patchNew_new_n348_);
  and eco173 (patchNew_new_n332_, g581, g4716);
  and eco174 (patchNew_new_n328_, g450, patchNew__not_GATE_24);
  not eco175 (patchNew__not_GATE_11, patchNew_new_n285_);
  and eco176 (patchNew_new_n272_, g610, g4767);
  and eco177 (patchNew_new_n318_, g4788, patchNew__not_GATE_20);
  and eco178 (patchNew_new_n273_, patchNew__not_GATE_6, patchNew_new_n272_);
  nor eco179 (patchNew_new_n351_, patchNew_new_n349_, patchNew_new_n350_);
  and eco180 (patchNew_new_n271_, g4814, g495);
  and eco181 (patchNew_new_n362_, g581, g4718);
  and eco182 (patchNew_new_n323_, g625, patchNew__not_GATE_22);
  and eco183 (patchNew_new_n304_, g4785, patchNew__not_GATE_16);
  nor eco184 (patchNew_new_n431_, patchNew_new_n429_, patchNew_new_n430_);
  and eco185 (patchNew_new_n432_, g4798, patchNew__not_GATE_54);
  and eco186 (patchNew_new_n262_, g4711, patchNew__not_GATE_0);
  not eco187 (patchNew__not_GATE_18, g4788);
  nor eco188 (patchNew_new_n285_, patchNew_new_n283_, patchNew_new_n284_);
  and eco189 (patchNew_new_n343_, g1068, g511_g4785_96);
  and eco190 (patchNew_new_n395_, g497, g4753);
  and eco191 (patchNew_new_n396_, patchNew__not_GATE_45, g4743);
  and eco192 (patchNew_new_n317_, g4785, g4727);
  and eco193 (patchNew_new_n310_, g4705, patchNew_new_n309_);
  nor eco194 (patchNew_new_n348_, g4788, g1035);
  and eco195 (patchNew_new_n268_, g4815, patchNew__not_GATE_4);
  not eco196 (patchNew__not_GATE_42, g4693);
  not eco197 (patchNew__not_GATE_9, patchNew_new_n275_);
  not eco198 (patchNew__not_GATE_48, g483);
  and eco199 (patchNew_new_n282_, g4813, patchNew__not_GATE_10);
  and eco200 (patchNew_new_n375_, g625, patchNew__not_GATE_39);
  not eco201 (patchNew__not_GATE_4, patchNew_new_n266_);
  nor eco202 (patchNew_new_n316_, g582, g730);
  nor eco203 (patchNew_new_n382_, g4791, patchNew_n321);
  and eco204 (patchNew_new_n384_, patchNew__not_GATE_42, g483);
  and eco205 (patchNew_new_n350_, g4701, patchNew_new_n309_);
  not eco206 (patchNew__not_GATE_7, patchNew_new_n274_);
  nor eco207 (patchNew_new_n344_, g4788, g4702_g4785_189);
  not eco208 (patchNew__not_GATE_16, patchNew_new_n303_);
  nor eco209 (patchNew_new_n307_, g4788, g648);
  nor eco210 (patchNew_new_n380_, patchNew_new_n375_, patchNew_new_n379_);
  and eco211 (patchNew_new_n280_, g609, g4746);
  not eco212 (patchNew__not_GATE_2, patchNew_new_n264_);
  nor eco213 (patchNew_new_n312_, patchNew_new_n308_, patchNew_new_n311_);
  not eco214 (patchNew__not_GATE_34, patchNew_new_n354_);
  not eco215 (patchNew__not_GATE_19, patchNew_new_n310_);
  nor eco216 (patchNew_new_n366_, g1015, patchNew_n373);
  and eco217 (patchNew_new_n264_, g4700, g4744);
  and eco218 (patchNew_new_n360_, g4785, patchNew__not_GATE_36);
  and eco219 (patchNew_new_n288_, g4814, g492);
  not eco220 (patchNew__not_GATE_32, patchNew_new_n346_);
  not eco221 (patchNew__not_GATE_50, g533);
  nor eco222 (patchNew_new_n321_, patchNew_new_n318_, patchNew_new_n320_);
  not eco223 (patchNew__not_GATE_91, g4785);
  and eco224 (patchNew_new_n541_, patchNew__not_GATE_92, g4709);
  not eco225 (patchNew__not_GATE_92, g4788);
  and eco226 (patchNew_new_n542_, g4785, patchNew__not_GATE_93);
  not eco227 (patchNew__not_GATE_93, patchNew_new_n541_);
  and eco228 (patchNew_new_n543_, g4741, g632);
  nor eco229 (patchNew_new_n544_, patchNew_new_n542_, patchNew_new_n543_);
  and eco230 (patchNew_new_n545_, g581, g4719);
  nor eco231 (patchNew_new_n546_, patchNew_new_n540_, patchNew_new_n545_);
  and eco232 (patchNew_new_n547_, patchNew__not_GATE_94, patchNew_new_n546_);
  and eco233 (patchNew_new_n548_, patchNew__not_GATE_95, patchNew_new_n547_);
  not eco234 (patchNew__not_GATE_94, patchNew_new_n544_);
  nor eco235 (patchNew_new_n429_, g510, patchNew_n1031);
  and eco236 (patchNew_new_n430_, g4683, g460);
  nor eco237 (patchNew_new_n393_, patchNew_new_n384_, patchNew_new_n392_);
  and eco238 (patchNew_new_n394_, g750, patchNew__not_GATE_44);
  and eco239 (patchNew_new_n397_, patchNew__not_GATE_46, g706);
  not eco240 (patchNew__not_GATE_46, g555);
  and eco241 (patchNew_new_n510_, patchNew__not_GATE_75, patchNew_new_n509_);
  not eco242 (patchNew__not_GATE_75, patchNew_new_n508_);
  nor eco243 (patchNew_new_n511_, patchNew_new_n505_, patchNew_new_n510_);
  and eco244 (patchNew_new_n512_, g4691, patchNew__not_GATE_76);
  nor eco245 (patchNew_new_n411_, patchNew_new_n407_, patchNew_new_n408_);
  nor eco246 (patchNew_new_n412_, patchNew_new_n409_, patchNew_new_n410_);
  and eco247 (patchNew_new_n489_, g581, g4710);
  and eco248 (patchNew_new_n414_, patchNew__not_GATE_48, patchNew_new_n413_);
  and eco249 (patchNew_new_n346_, patchNew__not_GATE_31, patchNew_new_n345_);
  not eco250 (patchNew__not_GATE_24, patchNew_new_n327_);
  and eco251 (patchNew_new_n330_, g542, patchNew__not_GATE_26);
  and eco252 (patchNew_new_n329_, patchNew__not_GATE_25, g4717);
  not eco253 (patchNew__not_GATE_8, patchNew_new_n273_);
  nor eco254 (patchNew_new_n476_, g491, g1123);
  and eco255 (patchNew_new_n477_, g706, patchNew__not_GATE_65);
  not eco256 (patchNew__not_GATE_65, g487);
  and eco257 (patchNew_new_n433_, g4680, patchNew__not_GATE_55);
  not eco258 (patchNew__not_GATE_54, patchNew_new_n431_);
  nor eco259 (patchNew_new_n466_, g1308, patchNew_new_n465_);
  nor eco260 (patchNew_new_n493_, patchNew_new_n491_, patchNew_new_n492_);
  not eco261 (patchNew__not_GATE_43, g483);
  nor eco262 (patchNew_new_n480_, patchNew_new_n477_, patchNew_new_n478_);
  and eco263 (patchNew_new_n481_, patchNew_new_n479_, patchNew_new_n480_);
  and eco264 (patchNew_new_n482_, patchNew__not_GATE_66, patchNew_new_n481_);
  and eco265 (patchNew_new_n445_, g4794, patchNew__not_GATE_58);
  not eco266 (patchNew__not_GATE_58, patchNew_new_n441_);
  and eco267 (patchNew_new_n424_, patchNew__not_GATE_52, patchNew_new_n423_);
  not eco268 (patchNew__not_GATE_45, g1123);
  and eco269 (patchNew_new_n340_, g630, g4735);
  and eco270 (patchNew_new_n284_, g4814, g4766);
  and eco271 (patchNew_new_n446_, g4680, patchNew_n348);
  and eco272 (patchNew_new_n447_, g4685, g643);
  not eco273 (patchNew__not_GATE_44, patchNew_new_n393_);
  and eco274 (patchNew_new_n354_, g576, g4740);
  and eco275 (patchNew_new_n472_, patchNew__not_GATE_64, patchNew_new_n393_);
  not eco276 (patchNew__not_GATE_64, g750);
  not eco277 (patchNew__not_GATE_23, patchNew_new_n321_);
  and eco278 (patchNew_new_n335_, g4785, g731);
  nor eco279 (patchNew_new_n305_, patchNew_new_n299_, patchNew_new_n300_);
  and eco280 (patchNew_new_n371_, g1340, patchNew_new_n364_);
  not eco281 (patchNew__not_GATE_56, g4798);
  not eco282 (patchNew__not_GATE_21, patchNew_new_n319_);
  and eco283 (patchNew_new_n289_, g4768, patchNew__not_GATE_12);
  and eco284 (patchNew_new_n410_, g1122, g4751);
  nor eco285 (patchNew_new_n387_, patchNew_n532, g476);
  and eco286 (patchNew_new_n386_, g1122, g4749);
  and eco287 (patchNew_new_n423_, g593, patchNew__not_GATE_51);
  not eco288 (patchNew__not_GATE_49, patchNew_new_n404_);
  not eco289 (patchNew__not_GATE_41, patchNew_new_n373_);
  nor eco290 (patchNew_new_n327_, g535, patchNew_new_n326_);
  and eco291 (patchNew_new_n462_, g685, patchNew__not_GATE_61);
  not eco292 (patchNew__not_GATE_61, patchNew_new_n415_);
  nor eco293 (patchNew_new_n296_, patchNew_new_n291_, patchNew_new_n295_);
  and eco294 (patchNew_new_n286_, g753, patchNew__not_GATE_11);
  nor eco295 (patchNew_new_n438_, patchNew_new_n436_, patchNew_new_n437_);
  nor eco296 (patchNew_new_n439_, g575, patchNew_new_n364_);
  and eco297 (patchNew_new_n294_, patchNew_new_n292_, patchNew_new_n293_);
  and eco298 (patchNew_new_n355_, g518, patchNew__not_GATE_34);
  and eco299 (patchNew_new_n283_, g4776, g705);
  and eco300 (patchNew_new_n385_, g4779, g471);
  and eco301 (patchNew_new_n368_, patchNew__not_GATE_38, patchNew_n244);
  and eco302 (patchNew_new_n263_, g4764, patchNew__not_GATE_1);
  nor eco303 (patchNew_new_n448_, patchNew_new_n446_, patchNew_new_n447_);
  nor eco304 (patchNew_new_n449_, g739, patchNew_new_n448_);
  and eco305 (patchNew_new_n314_, g581, g4715);
  and eco306 (patchNew_new_n363_, patchNew__not_GATE_37, patchNew_new_n362_);
  and eco307 (patchNew_new_n322_, g804, g4738);
  and eco308 (patchNew_new_n357_, g4788, patchNew__not_GATE_35);
  not eco309 (patchNew__not_GATE_31, patchNew_new_n343_);
  nor eco310 (patchNew_new_n389_, patchNew_new_n385_, patchNew_new_n386_);
  nor eco311 (patchNew_new_n390_, patchNew_new_n387_, patchNew_new_n388_);
  nor eco312 (patchNew_new_n339_, patchNew_new_n336_, patchNew_new_n338_);
  nor eco313 (patchNew_new_n490_, patchNew_new_n380_, patchNew_new_n489_);
  nor eco314 (patchNew_new_n491_, g445, patchNew_new_n490_);
  and eco315 (patchNew_new_n492_, g4681, g460);
  and eco316 (patchNew_new_n388_, g4769, g706);
  not eco317 (patchNew__not_GATE_13, g4814);
  and eco318 (patchNew_new_n290_, g4778, patchNew__not_GATE_13);
  and eco319 (patchNew_new_n292_, g4814, g478);
  and eco320 (patchNew_new_n421_, g569, patchNew__not_GATE_49);
  and eco321 (patchNew_new_n422_, patchNew__not_GATE_50, patchNew_n378);
  and eco322 (patchNew_new_n478_, g4775, g501);
  nor eco323 (patchNew_new_n479_, patchNew_new_n475_, patchNew_new_n476_);
  and eco324 (patchNew_new_n444_, g4797, patchNew__not_GATE_57);
  not eco325 (patchNew__not_GATE_57, patchNew_new_n423_);
  and eco326 (patchNew_new_n295_, g4813, patchNew__not_GATE_14);
  and eco327 (patchNew_new_n379_, g4785, patchNew__not_GATE_40);
  and eco328 (patchNew_new_n377_, g538, g4720);
  not eco329 (patchNew__not_GATE_40, patchNew_new_n378_);
  not eco330 (patchNew__not_GATE_12, patchNew_new_n288_);
  not eco331 (patchNew__not_GATE_66, g483);
  nor eco332 (patchNew_new_n483_, patchNew_new_n474_, patchNew_new_n482_);
  and eco333 (patchNew_new_n484_, g4691, patchNew__not_GATE_67);
  and eco334 (patchNew_new_n391_, patchNew_new_n389_, patchNew_new_n390_);
  and eco335 (patchNew_new_n417_, g4680, patchNew_n448);
  and eco336 (patchNew_new_n418_, g4674, g460);
  and eco337 (patchNew_new_n336_, g730, patchNew__not_GATE_28);
  not eco338 (patchNew__not_GATE_3, patchNew_new_n265_);
  and eco339 (patchNew_new_n265_, g4732, patchNew__not_GATE_2);
  not eco340 (patchNew__not_GATE_55, patchNew_n770);
  not eco341 (patchNew__not_GATE_5, patchNew_new_n263_);
  and eco342 (patchNew_new_n374_, g580, g4731);
  and eco343 (patchNew_new_n451_, g550, patchNew_new_n427_);
  nor eco344 (patchNew_new_n452_, patchNew_new_n428_, patchNew_new_n449_);
  and eco345 (patchNew_new_n313_, patchNew__not_GATE_19, patchNew_new_n312_);
  not eco346 (patchNew__not_GATE_33, g454);
  nor eco347 (patchNew_new_n372_, g1015, patchNew_new_n371_);
  and eco348 (patchNew_new_n408_, g4771, g706);
  nor eco349 (patchNew_new_n409_, patchNew_n532, g688);
  not eco350 (patchNew__not_GATE_14, patchNew_new_n294_);
  not eco351 (patchNew__not_GATE_29, patchNew_new_n337_);
  and eco352 (patchNew_new_n406_, patchNew__not_GATE_47, g483);
  not eco353 (patchNew__not_GATE_47, g4692);
  and eco354 (patchNew_new_n274_, g4814, g4757);
  not eco355 (patchNew__not_GATE_30, patchNew_new_n340_);
  and eco356 (patchNew_new_n401_, patchNew_new_n399_, patchNew_new_n400_);
  nor eco357 (patchNew_new_n352_, g448, patchNew_new_n351_);
  nor eco358 (patchNew_new_n436_, g4799, patchNew_new_n435_);
  and eco359 (patchNew_new_n437_, g4799, patchNew_new_n435_);
  and eco360 (patchNew_new_n319_, g4785, g4706);
  nor eco361 (patchNew_new_n291_, g4813, patchNew_new_n290_);
  and eco362 (patchNew_new_n338_, g4785, patchNew__not_GATE_29);
  and eco363 (patchNew_new_n426_, g4682, g624);
  nor eco364 (patchNew_new_n427_, patchNew_new_n425_, patchNew_new_n426_);
  and eco365 (patchNew_new_n293_, g4748, g4758);
  and eco366 (patchNew_new_n392_, patchNew__not_GATE_43, patchNew_new_n391_);
  not eco367 (patchNew__not_GATE_36, patchNew_new_n359_);
  not eco368 (patchNew__not_GATE_17, patchNew_new_n304_);
  and eco369 (patchNew_new_n266_, g4774, patchNew__not_GATE_3);
  nor eco370 (patchNew_new_n369_, g1015, patchNew_n1031);
  nor eco371 (patchNew_new_n453_, patchNew_new_n450_, patchNew_new_n451_);
  and eco372 (patchNew_new_n461_, patchNew_new_n457_, patchNew_new_n460_);
  nor eco373 (patchNew_new_n281_, patchNew_new_n279_, patchNew_new_n280_);
  and eco374 (patchNew_new_n471_, patchNew__not_GATE_63, patchNew_new_n465_);
  not eco375 (patchNew__not_GATE_63, g4808);
  and eco376 (patchNew_new_n407_, g4781, g471);
  and eco377 (patchNew_new_n378_, patchNew_new_n376_, patchNew_new_n377_);
  nor eco378 (patchNew_new_n364_, patchNew_new_n361_, patchNew_new_n363_);
  not eco379 (patchNew__not_GATE_20, patchNew_new_n317_);
  and eco380 (patchNew_new_n454_, patchNew_new_n452_, patchNew_new_n453_);
  not eco381 (patchNew__not_GATE_51, patchNew_new_n422_);
  and eco382 (patchNew_new_n496_, g505, g4677);
  and eco383 (patchNew_new_n405_, g4803, patchNew_new_n404_);
  nor eco384 (patchNew_new_n419_, patchNew_new_n417_, patchNew_new_n418_);
  nor eco385 (patchNew_new_n415_, patchNew_new_n406_, patchNew_new_n414_);
  and eco386 (patchNew_new_n416_, g686, patchNew_new_n415_);
  and eco387 (patchNew_new_n523_, patchNew__not_GATE_82, patchNew_new_n522_);
  not eco388 (patchNew__not_GATE_82, patchNew_new_n521_);
  nor eco389 (patchNew_new_n524_, patchNew_new_n520_, patchNew_new_n523_);
  nor eco390 (patchNew_new_n525_, patchNew_new_n394_, patchNew_new_n405_);
  nor eco391 (patchNew_new_n526_, patchNew_new_n416_, patchNew_new_n420_);
  not eco392 (patchNew__not_GATE_28, patchNew_new_n335_);
  and eco393 (patchNew_new_n499_, patchNew_new_n497_, patchNew__xnor_GATE_6);
  nor eco394 (patchNew_new_n500_, patchNew_new_n466_, patchNew_new_n483_);
  not eco395 (patchNew__not_GATE_6, patchNew_new_n271_);
  not eco396 (patchNew__not_GATE_35, patchNew_new_n356_);
  and eco397 (patchNew_new_n269_, g4787, patchNew__not_GATE_5);
  and eco398 (patchNew_new_n275_, g4813, patchNew__not_GATE_7);
  and eco399 (patchNew_new_n450_, patchNew__not_GATE_59, patchNew_new_n448_);
  not eco400 (patchNew__not_GATE_59, g4800);
  not eco401 (patchNew__not_GATE_53, patchNew_new_n427_);
  and eco402 (patchNew_new_n420_, g509, patchNew_new_n419_);
  and eco403 (patchNew_new_n434_, g4684, g665);
  nor eco404 (patchNew_new_n435_, patchNew_new_n433_, patchNew_new_n434_);
  not eco405 (patchNew__not_GATE_76, patchNew_new_n511_);
  and eco406 (patchNew_new_n513_, g4688, g687);
  nor eco407 (patchNew_new_n514_, patchNew_new_n512_, patchNew_new_n513_);
  and eco408 (patchNew_new_n460_, patchNew_new_n458_, patchNew_new_n459_);
  and eco409 (patchNew_new_n485_, g4694, g600);
  and eco410 (patchNew_new_n309_, g4785, patchNew__not_GATE_18);
  nor eco411 (patchNew_new_n463_, g483, patchNew_n747);
  and eco412 (patchNew_new_n464_, g4689, g483);
  nor eco413 (patchNew_new_n465_, patchNew_new_n463_, patchNew_new_n464_);
  nor eco414 (patchNew_new_n404_, patchNew_new_n402_, patchNew_new_n403_);
  not eco415 (patchNew__not_GATE_25, g730);
  nor eco416 (patchNew_new_n399_, patchNew_new_n395_, patchNew_new_n396_);
  nor eco417 (patchNew_new_n400_, patchNew_new_n397_, patchNew_new_n398_);
  nor eco418 (patchNew_new_n358_, patchNew_new_n355_, patchNew_new_n357_);
  and eco419 (patchNew_new_n277_, patchNew__not_GATE_8, patchNew_new_n276_);
  and eco420 (patchNew_new_n311_, g4788, g4726);
  and eco421 (patchNew_new_n504_, patchNew_new_n502_, patchNew_new_n503_);
  and eco422 (patchNew_new_n505_, g1122, g4750);
  and eco423 (patchNew_new_n506_, g4780, g501);
  and eco424 (patchNew_new_n507_, g4770, g706);
  xnor eco425 (patchNew__xnor_GATE_1, patchNew_n747, patchNew_new_n413_);
  xnor eco426 (patchNew__xnor_GATE_2, patchNew_new_n391_, patchNew_new_n401_);
  and eco427 (patchNew_new_n442_, g771, patchNew_new_n441_);
  and eco428 (patchNew_new_n443_, patchNew__not_GATE_56, patchNew_new_n431_);
  nor eco429 (patchNew_new_n373_, g633, g730);
  and eco430 (patchNew_new_n359_, g536, g4708);
  nor eco431 (patchNew_new_n467_, g553, patchNew_n1037);
  and eco432 (patchNew_new_n468_, g4695, g483);
  and eco433 (patchNew_new_n428_, g4796, patchNew__not_GATE_53);
  not eco434 (patchNew__not_GATE_26, patchNew_new_n329_);
  and eco435 (patchNew_new_n337_, g627, g4703);
  not eco436 (patchNew__not_GATE_22, patchNew_new_n322_);
  not eco437 (patchNew__not_GATE_37, patchNew_new_n361_);
  and eco438 (patchNew_new_n515_, g720, patchNew__not_GATE_77);
  not eco439 (patchNew__not_GATE_77, patchNew_new_n514_);
  and eco440 (patchNew_new_n516_, patchNew__not_GATE_78, patchNew_new_n514_);
  not eco441 (patchNew__not_GATE_78, g720);
  nor eco442 (patchNew_new_n486_, patchNew_new_n484_, patchNew_new_n485_);
  not eco443 (patchNew__not_GATE_67, patchNew_n477);
  nor eco444 (patchNew_new_n402_, g703, patchNew_new_n401_);
  and eco445 (patchNew_new_n403_, g4687, g483);
  and eco446 (patchNew_new_n457_, patchNew__not_GATE_60, patchNew_new_n456_);
  not eco447 (patchNew__not_GATE_60, patchNew_new_n444_);
  nor eco448 (patchNew_new_n469_, patchNew_new_n467_, patchNew_new_n468_);
  and eco449 (patchNew_new_n470_, patchNew__not_GATE_62, patchNew_new_n469_);
  not eco450 (patchNew__not_GATE_62, g4810);
  nor eco451 (patchNew_new_n473_, patchNew_new_n471_, patchNew_new_n472_);
  nor eco452 (patchNew_new_n474_, g904, patchNew_new_n469_);
  and eco453 (patchNew_new_n475_, g497, g4755);
  not eco454 (patchNew__not_GATE_38, g4791);
  and eco455 (patchNew_new_n519_, g461, patchNew__not_GATE_80);
  and eco456 (patchNew_new_n518_, patchNew__not_GATE_79, patchNew_n494);
  nor eco457 (patchNew_new_n522_, g509, patchNew_new_n419_);
  not eco458 (patchNew__not_GATE_79, g724);
  and eco459 (patchNew_new_n356_, g4785, g4729);
  and eco460 (patchNew_new_n458_, patchNew_new_n454_, patchNew_new_n455_);
  nor eco461 (patchNew_new_n459_, patchNew_new_n442_, patchNew_new_n445_);
  nor eco462 (patchNew_new_n527_, patchNew_new_n421_, patchNew_new_n462_);
  and eco463 (patchNew_new_n528_, patchNew_new_n526_, patchNew_new_n527_);
  and eco464 (patchNew_new_n529_, patchNew_new_n525_, patchNew_new_n528_);
  and eco465 (patchNew_new_n530_, patchNew__not_GATE_83, patchNew_new_n529_);
  not eco466 (patchNew__not_GATE_83, patchNew_new_n517_);
  and eco467 (patchNew_new_n508_, patchNew__not_GATE_74, g497);
  not eco468 (patchNew__not_GATE_74, g710);
  nor eco469 (patchNew_new_n509_, patchNew_new_n506_, patchNew_new_n507_);
  not eco470 (patchNew__not_GATE_80, patchNew_new_n518_);
  and eco471 (patchNew_new_n520_, g1332, patchNew_new_n519_);
  and eco472 (patchNew_new_n521_, g4802, patchNew__not_GATE_81);
  and eco473 (patchNew_new_n540_, patchNew__not_GATE_91, g4788);
  not eco474 (patchNew__not_GATE_81, patchNew_new_n519_);
  and eco475 (patchNew_new_n425_, g4680, patchNew_n244);
  not eco476 (patchNew__not_GATE_52, g4797);
  nor eco477 (patchNew_new_n361_, patchNew_new_n358_, patchNew_new_n360_);
  nor eco478 (patchNew_new_n345_, g1049, g1062);
  nor eco479 (patchNew_new_n455_, patchNew_new_n424_, patchNew_new_n432_);
  nor eco480 (patchNew_new_n456_, patchNew_new_n438_, patchNew_new_n443_);
  and eco481 (patchNew_new_n413_, patchNew_new_n411_, patchNew_new_n412_);
  and eco482 (patchNew_new_n502_, patchNew_new_n500_, patchNew__xnor_GATE_7);
  and eco483 (patchNew_new_n503_, patchNew__not_GATE_73, patchNew_new_n499_);
  not eco484 (patchNew__not_GATE_73, patchNew_new_n473_);
  and eco485 (patchNew_new_n531_, patchNew__not_GATE_84, patchNew_new_n530_);
  not eco486 (patchNew__not_GATE_84, patchNew_new_n524_);
  and eco487 (patchNew_new_n532_, patchNew__not_GATE_85, patchNew_new_n531_);
  not eco488 (patchNew__not_GATE_85, patchNew_new_n504_);
  not eco489 (patchNew__not_GATE_95, patchNew_new_n539_);
  nor eco490 (patchNew_new_n549_, g4790, patchNew__xnor_GATE_9);
  and eco491 (patchNew_new_n550_, g864, patchNew__not_GATE_96);
  not eco492 (patchNew__not_GATE_96, patchNew_new_n547_);
  and eco493 (patchNew_new_n551_, patchNew__not_GATE_97, patchNew_new_n550_);
  not eco494 (patchNew__not_GATE_97, patchNew_new_n549_);
  and eco495 (patchNew_new_n556_, patchNew_new_n481_, patchNew__xnor_GATE_8);
  nor eco496 (patchNew_new_n557_, patchNew_new_n481_, patchNew__xnor_GATE_8);
  nor eco497 (patchNew_new_n558_, patchNew_new_n556_, patchNew_new_n557_);
  not eco498 (patchNew__not_GATE_86, patchNew_new_n461_);
  and eco499 (patchNew_new_n534_, patchNew_new_n364_, patchNew__not_GATE_87);
  not eco500 (patchNew__not_GATE_87, patchNew_new_n490_);
  nor eco501 (patchNew_new_n535_, patchNew_n321, patchNew_new_n534_);
  and eco502 (patchNew_new_n539_, patchNew__not_GATE_90, patchNew__xnor_GATE_9);
  not eco503 (patchNew__not_GATE_90, g4790);
  and eco504 (patchNew_new_n619_, patchNew_n477, patchNew__not_GATE_123);
  not eco505 (patchNew__not_GATE_123, patchNew_new_n618_);
  and eco506 (patchNew_new_n620_, g4698, patchNew__not_GATE_124);
  not eco507 (patchNew__not_GATE_124, patchNew_new_n619_);
  and eco508 (patchNew_new_n621_, g569, patchNew_new_n620_);
  and eco509 (patchNew_new_n622_, patchNew_new_n617_, patchNew_new_n621_);
  and eco510 (patchNew_new_n623_, patchNew_new_n413_, patchNew_new_n622_);
  and eco511 (patchNew_new_n624_, g685, patchNew__not_GATE_125);
  not eco512 (patchNew__not_GATE_125, patchNew_new_n413_);
  and eco513 (patchNew_new_n625_, patchNew__not_GATE_126, patchNew_new_n413_);
  not eco514 (patchNew__not_GATE_126, g685);
  nor eco515 (patchNew_new_n626_, patchNew_new_n624_, patchNew_new_n625_);
  and eco516 (patchNew_new_n627_, patchNew__not_GATE_127, patchNew_new_n626_);
  not eco517 (patchNew__not_GATE_127, patchNew_new_n616_);
  and eco518 (patchNew_new_n628_, patchNew_new_n620_, patchNew__not_GATE_128);
  not eco519 (patchNew__not_GATE_128, patchNew_new_n627_);
  nor eco520 (patchNew_new_n629_, patchNew_new_n623_, patchNew_new_n628_);
  and eco521 (patchNew_new_n630_, g720, patchNew__not_GATE_129);
  not eco522 (patchNew__not_GATE_129, patchNew_new_n511_);
  and eco523 (patchNew_new_n631_, patchNew__not_GATE_130, patchNew_new_n511_);
  not eco524 (patchNew__not_GATE_130, g720);
  nor eco525 (patchNew_new_n632_, patchNew_new_n630_, patchNew_new_n631_);
  and eco526 (patchNew_new_n633_, patchNew__not_GATE_131, patchNew_new_n632_);
  not eco527 (patchNew__not_GATE_131, patchNew_new_n616_);
  and eco528 (patchNew_new_n634_, patchNew_new_n620_, patchNew_new_n633_);
  and eco529 (patchNew_new_n635_, patchNew__not_GATE_132, patchNew_new_n511_);
  not eco530 (patchNew__not_GATE_132, patchNew_new_n413_);
  and eco531 (patchNew_new_n636_, patchNew_new_n620_, patchNew_new_n635_);
  and eco532 (patchNew_new_n637_, patchNew_new_n634_, patchNew__not_GATE_133);
  not eco533 (patchNew__not_GATE_133, patchNew_new_n636_);
  nor eco534 (patchNew_new_n638_, patchNew_new_n629_, patchNew_new_n637_);
  and eco535 (patchNew_new_n639_, g1332, patchNew_new_n620_);
  and eco536 (patchNew_new_n640_, patchNew__not_GATE_134, patchNew_new_n639_);
  not eco537 (patchNew__not_GATE_134, patchNew_new_n616_);
  and eco538 (patchNew_new_n641_, patchNew__not_GATE_135, patchNew_new_n640_);
  not eco539 (patchNew__not_GATE_135, patchNew_n494);
  and eco540 (patchNew_new_n642_, patchNew_new_n614_, patchNew_new_n618_);
  and eco541 (patchNew_new_n643_, g509, patchNew__not_GATE_136);
  not eco542 (patchNew__not_GATE_136, patchNew_new_n642_);
  and eco543 (patchNew_new_n644_, g4676, patchNew__not_GATE_137);
  not eco544 (patchNew__not_GATE_137, patchNew_new_n643_);
  and eco545 (patchNew_new_n645_, g4676, patchNew__not_GATE_138);
  not eco546 (patchNew__not_GATE_138, patchNew_new_n616_);
  and eco547 (patchNew_new_n646_, patchNew_n448, patchNew__not_GATE_139);
  not eco548 (patchNew__not_GATE_139, patchNew_new_n645_);
  and eco549 (patchNew_new_n647_, patchNew__not_GATE_140, patchNew_new_n646_);
  not eco550 (patchNew__not_GATE_140, patchNew_new_n644_);
  and eco551 (patchNew_new_n648_, g739, patchNew__not_GATE_141);
  not eco552 (patchNew__not_GATE_141, patchNew_new_n642_);
  and eco553 (patchNew_new_n649_, g4676, patchNew__not_GATE_142);
  not eco554 (patchNew__not_GATE_142, patchNew_new_n648_);
  and eco555 (patchNew_new_n650_, patchNew_n348, patchNew__not_GATE_143);
  not eco556 (patchNew__not_GATE_143, patchNew_new_n645_);
  and eco557 (patchNew_new_n651_, patchNew_new_n649_, patchNew__not_GATE_144);
  not eco558 (patchNew__not_GATE_144, patchNew_new_n650_);
  and eco559 (patchNew_new_n652_, g658, patchNew__not_GATE_145);
  not eco560 (patchNew__not_GATE_145, patchNew_new_n642_);
  and eco561 (patchNew_new_n653_, g618, patchNew_new_n642_);
  nor eco562 (patchNew_new_n654_, patchNew_new_n652_, patchNew_new_n653_);
  and eco563 (patchNew_new_n655_, patchNew__not_GATE_146, patchNew_new_n654_);
  not eco564 (patchNew__not_GATE_146, patchNew_n1031);
  and eco565 (patchNew_new_n656_, patchNew_n1031, patchNew__not_GATE_147);
  not eco566 (patchNew__not_GATE_147, patchNew_new_n654_);
  and eco567 (patchNew_new_n657_, g813, patchNew__not_GATE_148);
  not eco568 (patchNew__not_GATE_148, patchNew_new_n642_);
  and eco569 (patchNew_new_n658_, g790, patchNew_new_n642_);
  nor eco570 (patchNew_new_n659_, patchNew_new_n657_, patchNew_new_n658_);
  nor eco571 (patchNew_new_n662_, patchNew_new_n655_, patchNew_new_n656_);
  and eco572 (patchNew_new_n664_, patchNew_new_n662_, patchNew__xnor_GATE_10);
  and eco573 (patchNew_new_n665_, patchNew_new_n651_, patchNew__not_GATE_151);
  not eco574 (patchNew__not_GATE_151, patchNew_new_n664_);
  and eco575 (patchNew_new_n666_, patchNew__not_GATE_152, patchNew_new_n650_);
  not eco576 (patchNew__not_GATE_152, patchNew_new_n649_);
  and eco577 (patchNew_new_n667_, patchNew_new_n656_, patchNew_new_n666_);
  nor eco578 (patchNew_new_n668_, patchNew_new_n665_, patchNew_new_n667_);
  and eco579 (patchNew_new_n669_, g4676, patchNew__not_GATE_153);
  not eco580 (patchNew__not_GATE_153, patchNew_new_n668_);
  and eco581 (patchNew_new_n670_, g4796, patchNew__not_GATE_154);
  not eco582 (patchNew__not_GATE_154, patchNew_new_n616_);
  and eco583 (patchNew_new_n671_, g4807, patchNew_new_n616_);
  nor eco584 (patchNew_new_n672_, patchNew_new_n670_, patchNew_new_n671_);
  and eco585 (patchNew_new_n673_, patchNew__not_GATE_155, patchNew_new_n672_);
  not eco586 (patchNew__not_GATE_155, patchNew_n244);
  and eco587 (patchNew_new_n674_, g4806, patchNew_new_n616_);
  and eco588 (patchNew_new_n675_, g4794, patchNew__not_GATE_156);
  not eco589 (patchNew__not_GATE_156, patchNew_new_n616_);
  and eco590 (patchNew_new_n676_, patchNew_n244, patchNew__not_GATE_157);
  not eco591 (patchNew__not_GATE_157, patchNew_new_n672_);
  nor eco592 (patchNew_new_n677_, patchNew_new_n674_, patchNew_new_n675_);
  and eco593 (patchNew_new_n678_, patchNew__not_GATE_158, patchNew_new_n677_);
  not eco594 (patchNew__not_GATE_158, patchNew_new_n676_);
  and eco595 (patchNew_new_n679_, patchNew_new_n364_, patchNew__not_GATE_159);
  not eco596 (patchNew__not_GATE_159, patchNew_new_n678_);
  nor eco597 (patchNew_new_n680_, patchNew_new_n673_, patchNew_new_n679_);
  and eco598 (patchNew_new_n681_, patchNew_new_n651_, patchNew__not_GATE_160);
  not eco599 (patchNew__not_GATE_160, patchNew_new_n680_);
  nor eco600 (patchNew_new_n682_, patchNew_new_n669_, patchNew_new_n681_);
  nor eco601 (patchNew_new_n683_, patchNew_new_n647_, patchNew_new_n682_);
  and eco602 (patchNew_new_n684_, patchNew__not_GATE_161, patchNew_new_n621_);
  not eco603 (patchNew__not_GATE_161, patchNew_new_n616_);
  and eco604 (patchNew_new_n685_, patchNew__not_GATE_162, patchNew_new_n620_);
  not eco605 (patchNew__not_GATE_162, patchNew_new_n617_);
  and eco606 (patchNew_new_n686_, patchNew__not_GATE_163, patchNew_new_n685_);
  not eco607 (patchNew__not_GATE_163, patchNew_new_n684_);
  nor eco608 (patchNew_new_n687_, patchNew_new_n622_, patchNew_new_n686_);
  and eco609 (patchNew_new_n688_, patchNew_new_n644_, patchNew__not_GATE_164);
  not eco610 (patchNew__not_GATE_164, patchNew_new_n646_);
  and eco611 (patchNew_new_n689_, patchNew_n494, patchNew__not_GATE_165);
  not eco612 (patchNew__not_GATE_165, patchNew_new_n616_);
  and eco613 (patchNew_new_n690_, patchNew_new_n620_, patchNew_new_n689_);
  and eco614 (patchNew_new_n691_, patchNew__not_GATE_166, patchNew_new_n690_);
  not eco615 (patchNew__not_GATE_166, patchNew_new_n639_);
  nor eco616 (patchNew_new_n692_, patchNew_new_n634_, patchNew_new_n688_);
  and eco617 (patchNew_new_n693_, patchNew__not_GATE_167, patchNew_new_n692_);
  not eco618 (patchNew__not_GATE_167, patchNew_new_n691_);
  and eco619 (patchNew_new_n694_, patchNew__not_GATE_168, patchNew_new_n693_);
  not eco620 (patchNew__not_GATE_168, patchNew_new_n641_);
  and eco621 (patchNew_new_n695_, patchNew_new_n687_, patchNew_new_n694_);
  and eco622 (patchNew_new_n696_, patchNew__not_GATE_169, patchNew_new_n695_);
  not eco623 (patchNew__not_GATE_169, patchNew_new_n683_);
  and eco624 (patchNew_new_n697_, patchNew__not_GATE_170, patchNew_new_n640_);
  not eco625 (patchNew__not_GATE_170, patchNew_new_n632_);
  nor eco626 (patchNew_new_n698_, patchNew_new_n690_, patchNew_new_n697_);
  and eco627 (patchNew_new_n699_, patchNew_new_n687_, patchNew_new_n698_);
  nor eco628 (patchNew_new_n700_, patchNew_new_n696_, patchNew_new_n699_);
  nor eco629 (patchNew_new_n701_, patchNew_new_n628_, patchNew_new_n700_);
  nor eco630 (patchNew_new_n703_, patchNew_new_n587_, patchNew_new_n591_);
  and eco631 (patchNew_new_n704_, patchNew_new_n587_, patchNew_new_n591_);
  nor eco632 (patchNew_new_n705_, patchNew_new_n703_, patchNew_new_n704_);
  and eco633 (patchNew_new_n706_, g581, g4715);
  and eco634 (patchNew_new_n707_, patchNew_new_n313_, patchNew__not_GATE_171);
  not eco635 (patchNew__not_GATE_171, patchNew_new_n706_);
  and eco636 (patchNew_new_n708_, patchNew__not_GATE_172, patchNew_new_n707_);
  not eco637 (patchNew__not_GATE_172, patchNew_n373);
  nor eco638 (patchNew_new_n709_, patchNew_n378, patchNew_new_n707_);
  nor eco639 (patchNew_new_n710_, patchNew_new_n708_, patchNew_new_n709_);
  and eco640 (patchNew_new_n714_, patchNew__not_GATE_175, patchNew__xnor_GATE_11);
  not eco641 (patchNew__not_GATE_175, patchNew_new_n605_);
  and eco642 (patchNew_new_n715_, patchNew_new_n605_, patchNew__not_GATE_176);
  not eco643 (patchNew__not_GATE_176, patchNew__xnor_GATE_11);
  nor eco644 (patchNew_new_n716_, g4697, patchNew_new_n714_);
  not eco645 (patchNew__not_GATE_177, patchNew_new_n716_);
  nor eco646 (patchNew_new_n718_, g923, g1240);
  and eco647 (patchNew_new_n719_, patchNew__not_GATE_178, patchNew_new_n718_);
  not eco648 (patchNew__not_GATE_178, patchNew_n1001);
  and eco649 (patchNew_new_n720_, g953, patchNew_n593);
  and eco650 (patchNew_new_n721_, patchNew_n835, patchNew_new_n720_);
  not eco651 (patchNew__not_GATE_179, patchNew_new_n719_);
  and eco652 (patchNew_new_n729_, g4669, g4671);
  and eco653 (patchNew_new_n730_, g4789, patchNew__not_GATE_182);
  not eco654 (patchNew__not_GATE_182, patchNew_new_n729_);
  not eco655 (patchNew__not_GATE_183, g4784);
  and eco656 (patchNew_new_n732_, g4807, g4808);
  not eco657 (patchNew__not_GATE_184, g4809);
  xnor eco658 (patchNew__xnor_GATE_0, g4811, patchNew_new_n481_);
  nand eco659 (patchNew_n532, g4813, g4814);
endmodule
