module top_eco(clk,\a[0] ,\a[1] ,\a[5] ,\b[0] ,\b[1] ,\b[2] ,\b[5] ,\op[0] ,\op[1] , n_523, n_568, wc1, n_522, n_525, n_534, n_569, n_570, n_571, wc8, n_590, n_594, n_596, n_558, n_545, n_531, n_554, n_521, n_739, n_718, n_551, n_593, n_676, n_539, n_780, wc52, wc54, wc55, wc58, overflow, greater,\y[6] ,\y[7] , less,\y[0] ,\y[1] ,\y[2] ,\y[3] ,\y[4] ,\y[5] , is_eq, n_854, n_855);
  input clk,\a[0] ,\a[1] ,\a[5] ;
  input \b[0] ,\b[1] ,\b[2] ,\b[5] ,\op[0] ;
  input \op[1] , n_523, n_568, wc1, n_522;
  input n_525, n_534, n_569, n_570, n_571;
  input wc8, n_590, n_594, n_596, n_558;
  input n_545, n_531, n_554, n_521, n_739;
  input n_718, n_551, n_593, n_676, n_539;
  input n_780, wc52, wc54, wc55, wc58;
  output overflow, greater,\y[6] ,\y[7] ;
  output less,\y[0] ,\y[1] ,\y[2] ,\y[3] ;
  output \y[4] ,\y[5] , is_eq, n_854, n_855;
  wire patchNew_add_28_29_n_21, patchNew_wc7, patchNew_n_113, patchNew_n_292;
  wire patchNew_n_295, patchNew_lt_44_17_n_37, patchNew_n_296, patchNew_wc0, patchNew_n_121;
  wire patchNew_n_298, patchNew_n_301, patchNew_sub_33_29_n_54, patchNew_lt_44_17_n_71, patchNew_n_276;
  wire patchNew_n_241, patchNew_wc3, patchNew_n_110, patchNew_wc4, patchNew_n_510;
  wire patchNew_n_505, patchNew_wc5, patchNew_temp_y5, patchNew_temp_y0, patchNew_n_506;
  wire patchNew_wc6, patchNew_n_495, patchNew_n_496, patchNew_n_508, patchNew_n_426;
  wire patchNew_n_258, patchNew_n_438, patchNew_n_109, patchNew_n_242, patchNew_n_509;
  wire patchNew_wc8, patchNew_n_511, patchNew_wc9, patchNew_temp_y1, patchNew_temp_y4;
  wire patchNew_n_283, patchNew_wc10, patchNew_n_513, patchNew_wc11, patchNew_temp_y2;
  wire patchNew_temp_y3, patchNew_n_514, patchNew_wc12, patchNew_wc13, patchNew_n_489;
  wire patchNew_n_483, patchNew_n_484, patchNew_n_287, patchNew_n_490, patchNew_n_477;
  wire patchNew_n_478, patchNew_n_253, patchNew_wc14, patchNew_wc16, patchNew_wc15;
  wire patchNew_n_281, patchNew_n_456, patchNew_n_252, patchNew_n_278, patchNew_n_457;
  wire patchNew_n_472, patchNew_wc17, patchNew_n_450, patchNew_n_521, patchNew_sub_33_29_n_67;
  wire patchNew_n_522, patchNew_add_28_29_n_60, patchNew_n_451, patchNew_n_524, patchNew_wc18;
  wire patchNew_wc20, patchNew_n_525, patchNew_wc19, patchNew_n_462, patchNew_n_463;
  wire patchNew_n_358, patchNew_n_468, patchNew_n_469, patchNew_wc21, patchNew_n_254;
  wire patchNew_n_257, patchNew_lt_44_17_n_36, patchNew_n_418, patchNew_gt_43_12_n_36, patchNew_lt_44_17_n_88;
  wire patchNew_n_442, patchNew_wc22, patchNew_n_427, patchNew_n_306, patchNew_n_360;
  wire patchNew_wc44, patchNew_n_362, patchNew_wc43, patchNew_n_439, patchNew_n_285;
  wire patchNew_n_445, patchNew_n_255, patchNew_wc23, patchNew_lt_44_17_n_44, patchNew_n_421;
  wire patchNew_n_294, patchNew_add_28_29_n_47, patchNew_lt_44_17_n_87, patchNew_wc25, patchNew_add_28_29_n_50;
  wire patchNew_n_527, patchNew_n_289, patchNew_n_300, patchNew_gt_43_12_n_87, patchNew_n_528;
  wire patchNew_wc26, patchNew_add_28_29_n_56, patchNew_wc27, patchNew_n_530, patchNew_n_432;
  wire patchNew_n_433, patchNew_n_529, patchNew_wc28, patchNew_n_533, patchNew_n_531;
  wire patchNew_n_532, patchNew_sub_33_29_n_63, patchNew_n_534, patchNew_n_402, patchNew_n_397;
  wire patchNew_n_244, patchNew_lt_44_17_n_66, patchNew_n_412, patchNew_gt_43_12_n_66, patchNew_n_403;
  wire patchNew_n_394, patchNew_n_299, patchNew_n_409, patchNew_n_406, patchNew_sub_33_29_n_48;
  wire patchNew_gt_43_12_n_65, patchNew_n_293, patchNew_lt_44_17_n_65, patchNew_add_28_29_n_41, patchNew_n_260;
  wire patchNew_n_290, patchNew_n_536, patchNew_n_535, patchNew_n_537, patchNew_wc30;
  wire patchNew_n_259, patchNew_n_538, patchNew_wc31, patchNew_n_539, patchNew_wc32;
  wire patchNew_n_243, patchNew_sub_33_29_n_32, patchNew_sub_33_29_n_60, patchNew_n_540, patchNew_n_541;
  wire patchNew_n_542, patchNew_wc34, patchNew_add_28_29_n_53, patchNew_n_318, patchNew_wc35;
  wire patchNew_n_325, patchNew_n_502, patchNew_n_286, patchNew_n_499, patchNew_n_369;
  wire patchNew_n_370, patchNew_n_381, patchNew_n_382, patchNew_n_390, patchNew_n_391;
  wire patchNew_n_375, patchNew_n_376, patchNew_n_280, patchNew_wc36, patchNew_n_359;
  wire patchNew_wc37, patchNew_n_284, patchNew_n_249, patchNew_n_297, patchNew_gt_43_12_n_34;
  wire patchNew_n_282, patchNew_n_288, patchNew_n_389, patchNew_n_543, patchNew_n_354;
  wire patchNew_n_355, patchNew_n_330, patchNew_n_331, patchNew_n_342, patchNew_n_343;
  wire patchNew_n_348, patchNew_n_349, patchNew_n_368, patchNew_wc39, patchNew_n_363;
  wire patchNew_wc40, patchNew_n_544, patchNew_wc41, patchNew_n_364, patchNew_wc42;
  wire patchNew_n_361, patchNew_n_336, patchNew_n_337, patchNew_wc45, patchNew_add_28_29_n_51;
  wire patchNew_wc46, patchNew_n_312, patchNew_lt_44_17_n_68, patchNew_wc51, patchNew_wc53;
  wire patchNew_wc52, patchNew_wc54, patchNew_wc57, patchNew_wc55, patchNew_wc56;
  wire patchNew_n_34, patchNew_n_346, patchNew_n_347, patchNew_n_308, patchNew_n_307;
  wire patchNew_n_27, patchNew_n_24, patchNew_add_28_29_n_45, patchNew_n_323, patchNew_n_317;
  wire patchNew_n_320, patchNew_wc58, patchNew_n_332, patchNew_n_262, patchNew_add_28_29_n_44;
  wire patchNew_n_415, patchNew_wc65, patchNew_wc66, patchNew_wc67;
  and eco1 (\y[0] , patchNew_temp_y0, patchNew_wc53);
  and eco2 (\y[1] , patchNew_temp_y1, patchNew_wc52);
  and eco3 (\y[2] , patchNew_wc54, patchNew_temp_y2);
  and eco4 (\y[3] , patchNew_wc55, patchNew_temp_y3);
  and eco5 (\y[4] , patchNew_wc56, patchNew_temp_y4);
  and eco6 (\y[5] , patchNew_wc57, patchNew_temp_y5);
  and eco7 (is_eq, patchNew_gt_43_12_n_36, patchNew_lt_44_17_n_36);
  or eco8 (n_854, patchNew_wc3, patchNew_n_110);
  or eco9 (n_855, patchNew_n_241, patchNew_wc4);
  nand eco10 (patchNew_add_28_29_n_21,\a[0] , patchNew_n_113);
  assign overflow = \y[7] ;
  not eco12 (greater, patchNew_gt_43_12_n_36);
  nor eco13 (\y[6] , patchNew_n_472, patchNew_n_358);
  not eco14 (\y[7] , patchNew_n_358);
  and eco15 (less, patchNew_gt_43_12_n_36, patchNew_wc51);
  not eco16 (patchNew_wc7, patchNew_n_242);
  nand eco17 (patchNew_n_113, patchNew_n_306, patchNew_n_360);
  nand eco18 (patchNew_n_292, patchNew_n_113, patchNew_lt_44_17_n_37);
  or eco19 (patchNew_n_295, patchNew_wc0,\a[1] );
  not eco20 (patchNew_lt_44_17_n_37,\a[0] );
  or eco21 (patchNew_n_296, patchNew_n_121,\a[1] );
  not eco22 (patchNew_wc0, patchNew_n_121);
  nand eco23 (patchNew_n_121, patchNew_n_361, patchNew_n_362);
  or eco24 (patchNew_n_298, patchNew_n_113, wc52);
  nand eco25 (patchNew_n_301, patchNew_sub_33_29_n_54, patchNew_lt_44_17_n_71);
  nand eco26 (patchNew_sub_33_29_n_54, patchNew_lt_44_17_n_66, patchNew_n_412);
  not eco27 (patchNew_lt_44_17_n_71, patchNew_n_262);
  nand eco28 (patchNew_n_241, patchNew_n_505, patchNew_n_506);
  not eco29 (patchNew_wc3, patchNew_n_241);
  nand eco30 (patchNew_n_110, patchNew_n_508, patchNew_n_509);
  not eco31 (patchNew_wc4, patchNew_n_110);
  or eco32 (patchNew_n_510, patchNew_wc9, patchNew_temp_y1);
  or eco33 (patchNew_n_505, patchNew_wc5, patchNew_temp_y5);
  not eco34 (patchNew_wc5, patchNew_temp_y0);
  nand eco35 (patchNew_temp_y5, patchNew_n_495, patchNew_n_496);
  nand eco36 (patchNew_temp_y0, patchNew_n_390, patchNew_n_391);
  or eco37 (patchNew_n_506, patchNew_temp_y0, patchNew_wc6);
  not eco38 (patchNew_wc6, patchNew_temp_y5);
  or eco39 (patchNew_n_495,\op[1] , patchNew_wc13);
  nand eco40 (patchNew_n_496, patchNew_n_284,\op[1] );
  or eco41 (patchNew_n_508, patchNew_wc7, patchNew_n_109);
  nand eco42 (patchNew_n_426, patchNew_add_28_29_n_47, patchNew_add_28_29_n_50);
  nand eco43 (patchNew_n_258, patchNew_n_533, patchNew_n_534);
  or eco44 (patchNew_n_438,\op[1] , patchNew_wc25);
  nand eco45 (patchNew_n_109, patchNew_n_513, patchNew_n_514);
  nand eco46 (patchNew_n_242, patchNew_n_510, patchNew_n_511);
  or eco47 (patchNew_n_509, patchNew_n_242, patchNew_wc8);
  not eco48 (patchNew_wc8, patchNew_n_109);
  or eco49 (patchNew_n_511, patchNew_temp_y4, patchNew_wc10);
  not eco50 (patchNew_wc9, patchNew_temp_y4);
  nand eco51 (patchNew_temp_y1, patchNew_n_438, patchNew_n_439);
  nand eco52 (patchNew_temp_y4, patchNew_n_489, patchNew_n_490);
  nand eco53 (patchNew_n_283, patchNew_n_477, patchNew_n_478);
  not eco54 (patchNew_wc10, patchNew_temp_y1);
  or eco55 (patchNew_n_513, patchNew_wc11, patchNew_temp_y2);
  not eco56 (patchNew_wc11, patchNew_temp_y3);
  nand eco57 (patchNew_temp_y2, patchNew_n_462, patchNew_n_463);
  nand eco58 (patchNew_temp_y3, patchNew_n_483, patchNew_n_484);
  or eco59 (patchNew_n_514, patchNew_temp_y3, patchNew_wc12);
  not eco60 (patchNew_wc12, patchNew_temp_y2);
  not eco61 (patchNew_wc13, patchNew_n_283);
  or eco62 (patchNew_n_489,\op[1] , patchNew_wc14);
  or eco63 (patchNew_n_483,\op[1] , patchNew_wc15);
  nand eco64 (patchNew_n_484, patchNew_n_282,\op[1] );
  nand eco65 (patchNew_n_287, patchNew_n_456, patchNew_n_457);
  nand eco66 (patchNew_n_490, patchNew_n_288,\op[1] );
  or eco67 (patchNew_n_477, patchNew_wc16,\op[0] );
  nand eco68 (patchNew_n_478, patchNew_n_253,\op[0] );
  nand eco69 (patchNew_n_253, patchNew_n_521, patchNew_n_522);
  not eco70 (patchNew_wc14, patchNew_n_287);
  not eco71 (patchNew_wc16, patchNew_n_252);
  not eco72 (patchNew_wc15, patchNew_n_281);
  nand eco73 (patchNew_n_281, patchNew_n_450, patchNew_n_451);
  or eco74 (patchNew_n_456, patchNew_wc20,\op[0] );
  nand eco75 (patchNew_n_252, patchNew_n_524, patchNew_n_525);
  or eco76 (patchNew_n_278, patchNew_wc22, patchNew_n_427);
  nand eco77 (patchNew_n_457, patchNew_n_255,\op[0] );
  or eco78 (patchNew_n_472, patchNew_wc17,\op[1] );
  not eco79 (patchNew_wc17, patchNew_n_278);
  or eco80 (patchNew_n_450, patchNew_wc21,\op[0] );
  nand eco81 (patchNew_n_521, patchNew_sub_33_29_n_67, n_558);
  nand eco82 (patchNew_sub_33_29_n_67, n_521, patchNew_n_418);
  or eco83 (patchNew_n_522, patchNew_sub_33_29_n_67, n_558);
  nand eco84 (patchNew_add_28_29_n_60, n_739, patchNew_n_421);
  nand eco85 (patchNew_n_451, patchNew_n_258,\op[0] );
  or eco86 (patchNew_n_524, patchNew_wc18, n_558);
  not eco87 (patchNew_wc18, patchNew_add_28_29_n_60);
  not eco88 (patchNew_wc20, patchNew_n_254);
  or eco89 (patchNew_n_525, patchNew_add_28_29_n_60, patchNew_wc19);
  not eco90 (patchNew_wc19, n_558);
  or eco91 (patchNew_n_462,\op[1] , patchNew_wc23);
  nand eco92 (patchNew_n_463, patchNew_n_286,\op[1] );
  or eco93 (patchNew_n_358, patchNew_n_468, patchNew_n_469);
  or eco94 (patchNew_n_468, patchNew_wc65,\op[1] );
  nand eco95 (patchNew_n_469,\op[0] , patchNew_lt_44_17_n_68);
  not eco96 (patchNew_wc21, patchNew_n_257);
  nand eco97 (patchNew_n_254, patchNew_n_529, patchNew_n_530);
  nand eco98 (patchNew_n_257, patchNew_n_527, patchNew_n_528);
  nand eco99 (patchNew_lt_44_17_n_36, patchNew_lt_44_17_n_88, patchNew_n_442);
  nand eco100 (patchNew_n_418, patchNew_sub_33_29_n_54, n_522);
  nand eco101 (patchNew_gt_43_12_n_36, n_593, patchNew_n_445);
  nand eco102 (patchNew_lt_44_17_n_88, patchNew_n_346, patchNew_n_347);
  nand eco103 (patchNew_n_442, patchNew_n_294, patchNew_lt_44_17_n_87);
  not eco104 (patchNew_wc22, patchNew_n_426);
  or eco105 (patchNew_n_427, patchNew_wc45,\op[0] );
  or eco106 (patchNew_n_306, wc8, clk);
  nand eco107 (patchNew_n_360,\b[0] , clk);
  not eco108 (patchNew_wc44,\a[0] );
  nand eco109 (patchNew_n_362,\b[1] , clk);
  not eco110 (patchNew_wc43, n_539);
  nand eco111 (patchNew_n_439, patchNew_n_290,\op[1] );
  nand eco112 (patchNew_n_285, patchNew_n_432, patchNew_n_433);
  nand eco113 (patchNew_n_445, patchNew_n_300, patchNew_gt_43_12_n_87);
  nand eco114 (patchNew_n_255, patchNew_n_531, patchNew_n_532);
  not eco115 (patchNew_wc23, patchNew_n_285);
  nand eco116 (patchNew_n_421, patchNew_add_28_29_n_47, n_590);
  nand eco117 (patchNew_n_294, patchNew_lt_44_17_n_66, patchNew_n_406);
  nand eco118 (patchNew_add_28_29_n_47, patchNew_add_28_29_n_45, patchNew_n_415);
  nor eco119 (patchNew_lt_44_17_n_87, patchNew_n_262, patchNew_n_307);
  not eco120 (patchNew_wc25, patchNew_n_289);
  and eco121 (patchNew_add_28_29_n_50, patchNew_n_312, n_590);
  or eco122 (patchNew_n_527, patchNew_wc26, n_554);
  nand eco123 (patchNew_n_289, patchNew_n_402, patchNew_n_403);
  nand eco124 (patchNew_n_300, patchNew_gt_43_12_n_66, patchNew_n_409);
  nor eco125 (patchNew_gt_43_12_n_87, patchNew_n_332, patchNew_n_308);
  or eco126 (patchNew_n_528, patchNew_add_28_29_n_56, patchNew_wc27);
  not eco127 (patchNew_wc26, patchNew_add_28_29_n_56);
  nand eco128 (patchNew_add_28_29_n_56, n_676, patchNew_n_397);
  not eco129 (patchNew_wc27, n_554);
  or eco130 (patchNew_n_530, patchNew_add_28_29_n_47, patchNew_wc66);
  or eco131 (patchNew_n_432, patchNew_wc67,\op[0] );
  nand eco132 (patchNew_n_433, patchNew_n_244,\op[0] );
  or eco133 (patchNew_n_529, patchNew_wc28, n_545);
  not eco134 (patchNew_wc28, patchNew_add_28_29_n_47);
  nand eco135 (patchNew_n_533, patchNew_sub_33_29_n_63, n_554);
  nand eco136 (patchNew_n_531, patchNew_sub_33_29_n_54, n_545);
  or eco137 (patchNew_n_532, patchNew_sub_33_29_n_54, n_545);
  nand eco138 (patchNew_sub_33_29_n_63, patchNew_lt_44_17_n_44, patchNew_n_394);
  or eco139 (patchNew_n_534, patchNew_sub_33_29_n_63, n_554);
  or eco140 (patchNew_n_402, patchNew_wc30,\op[0] );
  nand eco141 (patchNew_n_397, patchNew_add_28_29_n_41, n_596);
  nand eco142 (patchNew_n_244, patchNew_n_535, patchNew_n_536);
  nand eco143 (patchNew_lt_44_17_n_66, patchNew_n_24, n_523);
  nand eco144 (patchNew_n_412, patchNew_sub_33_29_n_48, patchNew_lt_44_17_n_65);
  nand eco145 (patchNew_gt_43_12_n_66, patchNew_n_27, n_531);
  nand eco146 (patchNew_n_403, patchNew_n_260,\op[0] );
  nand eco147 (patchNew_n_394, patchNew_sub_33_29_n_48, n_525);
  nand eco148 (patchNew_n_299, patchNew_n_381, patchNew_n_382);
  nand eco149 (patchNew_n_409, patchNew_n_299, patchNew_gt_43_12_n_65);
  nand eco150 (patchNew_n_406, patchNew_n_293, patchNew_lt_44_17_n_65);
  nand eco151 (patchNew_sub_33_29_n_48, patchNew_n_318, patchNew_n_499);
  not eco152 (patchNew_gt_43_12_n_65, patchNew_n_24);
  nand eco153 (patchNew_n_293, patchNew_n_375, patchNew_n_376);
  not eco154 (patchNew_lt_44_17_n_65, patchNew_n_27);
  nand eco155 (patchNew_add_28_29_n_41, patchNew_n_325, patchNew_n_502);
  nand eco156 (patchNew_n_260, patchNew_n_539, patchNew_n_540);
  nand eco157 (patchNew_n_290, patchNew_n_369, patchNew_n_370);
  or eco158 (patchNew_n_536, patchNew_sub_33_29_n_48, n_551);
  nand eco159 (patchNew_n_535, patchNew_sub_33_29_n_48, n_551);
  or eco160 (patchNew_n_537, patchNew_wc31, n_551);
  not eco161 (patchNew_wc30, patchNew_n_259);
  nand eco162 (patchNew_n_259, patchNew_n_541, patchNew_n_542);
  or eco163 (patchNew_n_538, patchNew_add_28_29_n_41, patchNew_wc32);
  not eco164 (patchNew_wc31, patchNew_add_28_29_n_41);
  nand eco165 (patchNew_n_539, patchNew_sub_33_29_n_32, patchNew_sub_33_29_n_60);
  not eco166 (patchNew_wc32, n_551);
  nand eco167 (patchNew_n_243, patchNew_n_537, patchNew_n_538);
  nand eco168 (patchNew_sub_33_29_n_32, patchNew_lt_44_17_n_37, patchNew_n_113);
  nand eco169 (patchNew_sub_33_29_n_60, patchNew_n_318, patchNew_n_295);
  or eco170 (patchNew_n_540, patchNew_sub_33_29_n_32, patchNew_sub_33_29_n_60);
  or eco171 (patchNew_n_541, patchNew_wc34, patchNew_add_28_29_n_53);
  or eco172 (patchNew_n_542, patchNew_add_28_29_n_21, patchNew_wc35);
  not eco173 (patchNew_wc34, patchNew_add_28_29_n_21);
  nand eco174 (patchNew_add_28_29_n_53, patchNew_n_296, patchNew_n_325);
  or eco175 (patchNew_n_318, patchNew_n_121, wc54);
  not eco176 (patchNew_wc35, patchNew_add_28_29_n_53);
  nand eco177 (patchNew_n_325, patchNew_n_121,\a[1] );
  or eco178 (patchNew_n_502, patchNew_wc36, patchNew_add_28_29_n_21);
  nand eco179 (patchNew_n_286, patchNew_n_348, patchNew_n_349);
  nand eco180 (patchNew_n_499, patchNew_n_295, patchNew_sub_33_29_n_32);
  or eco181 (patchNew_n_369, patchNew_n_368, patchNew_wc39);
  nand eco182 (patchNew_n_370, patchNew_n_249,\op[0] );
  nand eco183 (patchNew_n_381, patchNew_n_298, patchNew_gt_43_12_n_34);
  nand eco184 (patchNew_n_382, patchNew_n_297, patchNew_n_121);
  or eco185 (patchNew_n_390, patchNew_n_389, patchNew_n_113);
  nand eco186 (patchNew_n_391, patchNew_n_280, patchNew_n_113);
  nand eco187 (patchNew_n_375, patchNew_n_292,\a[1] );
  or eco188 (patchNew_n_376, patchNew_wc37, patchNew_n_121);
  nand eco189 (patchNew_n_280, patchNew_n_330, patchNew_n_331);
  not eco190 (patchNew_wc36, patchNew_n_296);
  or eco191 (patchNew_n_359, patchNew_n_363, patchNew_wc42);
  not eco192 (patchNew_wc37, patchNew_n_359);
  nand eco193 (patchNew_n_284, patchNew_n_342, patchNew_n_343);
  nand eco194 (patchNew_n_249, patchNew_n_543, patchNew_n_544);
  or eco195 (patchNew_n_297, patchNew_n_364, patchNew_n_113);
  not eco196 (patchNew_gt_43_12_n_34,\a[1] );
  nand eco197 (patchNew_n_282, patchNew_n_336, patchNew_n_337);
  nand eco198 (patchNew_n_288, patchNew_n_354, patchNew_n_355);
  nand eco199 (patchNew_n_389,\a[0] , n_539);
  or eco200 (patchNew_n_543, patchNew_wc40, patchNew_n_121);
  or eco201 (patchNew_n_354,\op[0] , n_739);
  nand eco202 (patchNew_n_355, n_545,\op[0] );
  or eco203 (patchNew_n_330, n_539, patchNew_wc44);
  or eco204 (patchNew_n_331, patchNew_wc43,\a[0] );
  or eco205 (patchNew_n_342,\op[0] , n_780);
  nand eco206 (patchNew_n_343, n_558,\op[0] );
  or eco207 (patchNew_n_348,\op[0] , n_676);
  nand eco208 (patchNew_n_349, n_551,\op[0] );
  or eco209 (patchNew_n_368, patchNew_wc46,\op[0] );
  not eco210 (patchNew_wc39, patchNew_n_121);
  or eco211 (patchNew_n_363,\a[1] ,\a[0] );
  not eco212 (patchNew_wc40,\a[1] );
  or eco213 (patchNew_n_544,\a[1] , patchNew_wc41);
  not eco214 (patchNew_wc41, patchNew_n_121);
  nand eco215 (patchNew_n_364,\a[1] ,\a[0] );
  not eco216 (patchNew_wc42, patchNew_n_113);
  or eco217 (patchNew_n_361, wc1, clk);
  or eco218 (patchNew_n_336,\op[0] , n_718);
  nand eco219 (patchNew_n_337, n_554,\op[0] );
  not eco220 (patchNew_wc45, patchNew_add_28_29_n_51);
  nand eco221 (patchNew_add_28_29_n_51, patchNew_n_312, patchNew_n_320);
  not eco222 (patchNew_wc46,\a[1] );
  or eco223 (patchNew_n_312,\b[5] ,\a[5] );
  not eco224 (patchNew_lt_44_17_n_68, patchNew_n_34);
  not eco225 (patchNew_wc51, patchNew_lt_44_17_n_36);
  not eco226 (patchNew_wc53, patchNew_n_358);
  not eco227 (patchNew_wc52, patchNew_n_358);
  not eco228 (patchNew_wc54, patchNew_n_358);
  not eco229 (patchNew_wc57, patchNew_n_358);
  not eco230 (patchNew_wc55, patchNew_n_358);
  not eco231 (patchNew_wc56, patchNew_n_358);
  nand eco232 (patchNew_n_34, patchNew_n_317, patchNew_n_276);
  or eco233 (patchNew_n_346, patchNew_n_34, patchNew_n_308);
  nand eco234 (patchNew_n_347, n_569, patchNew_n_307);
  nand eco235 (patchNew_n_27, n_523, n_525);
  nand eco236 (patchNew_n_24, n_531, patchNew_lt_44_17_n_44);
  nand eco237 (patchNew_add_28_29_n_45, n_594, patchNew_n_323);
  nand eco238 (patchNew_n_323, n_676, n_718);
  or eco239 (patchNew_n_317, n_521, patchNew_wc58);
  nand eco240 (patchNew_n_320, n_739, n_780);
  not eco241 (patchNew_wc58, n_534);
  nand eco242 (patchNew_n_332, n_521, patchNew_n_276);
  nand eco243 (patchNew_n_262, n_522, n_534);
  and eco244 (patchNew_add_28_29_n_44, n_594, n_596);
  nand eco245 (patchNew_n_415, patchNew_add_28_29_n_41, patchNew_add_28_29_n_44);
  not eco246 (patchNew_wc65, patchNew_n_301);
  not eco247 (patchNew_wc66, n_545);
  not eco248 (patchNew_wc67, patchNew_n_243);
  nand eco249 (patchNew_n_307, n_568, n_570);
  nand eco250 (patchNew_n_308, n_569, n_571);
  or eco251 (patchNew_lt_44_17_n_44, wc55,\b[2] );
  or eco252 (patchNew_n_276,\b[5] , wc58);
endmodule
