module top(clk, oe, a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], b[0], b[1], b[2], b[3], b[4], b[5], b[6], b[7], op[0], op[1], y[0], y[1], y[2], y[3], y[4], y[5], y[6], y[7], parity, overflow, greater, is_eq, less);
  input clk, oe, a[0], a[1], a[2], a[3];
  input a[4], a[5], a[6], a[7], b[0], b[1];
  input b[2], b[3], b[4], b[5], b[6], b[7];
  input op[0], op[1];
  output y[0], y[1], y[2], y[3], y[4], y[5];
  output y[6], y[7], parity, overflow, greater, is_eq;
  output less;
  or eco1 (n_506, b[1], wc0);
  nand eco2 (parity, n_803, n_804);
  assign overflow = y[7];
  and eco4 (y[0], n_495, patchNew_wc66);
  and eco5 (greater, wc70, n_517);
  and eco6 (y[1], n_508, patchNew_wc63);
  and eco7 (y[2], n_480, patchNew_wc68);
  and eco8 (y[3], n_492, patchNew_wc67);
  and eco9 (y[4], n_488, patchNew_wc65);
  and eco10 (y[5], patchNew_wc69, n_504);
  assign y[6] = y[7];
  not eco12 (y[7], patchNew_n_69);
  nor eco13 (is_eq, n_517, n_520);
  and eco14 (less, wc69, n_520);
  nand eco15 (n_496, n_845, n_846);
  or eco16 (n_505, wc, a[1]);
  not eco17 (wc, b[1]);
  or eco18 (n_474, wc2, a[2]);
  not eco19 (wc0, a[1]);
  or eco20 (n_473, b[2], wc1);
  not eco21 (wc1, a[2]);
  or eco22 (n_481, b[4], wc3);
  not eco23 (wc2, b[2]);
  or eco24 (n_482, wc4, a[4]);
  not eco25 (wc3, a[4]);
  or eco26 (n_489, wc5, a[3]);
  not eco27 (wc4, b[4]);
  or eco28 (n_490, b[3], wc6);
  not eco29 (wc5, b[3]);
  not eco30 (wc6, a[3]);
  nand eco31 (n_537, n_473, n_506);
  or eco32 (n_515, b[5], wc7);
  not eco33 (wc7, a[5]);
  nand eco34 (n_539, n_474, n_505);
  or eco35 (n_542, n_483, a[3]);
  or eco36 (n_541, a[2], n_475);
  nand eco37 (n_475, n_851, n_852);
  or eco38 (n_543, n_477, a[1]);
  nand eco39 (n_483, n_837, n_838);
  nand eco40 (n_477, n_849, n_850);
  or eco41 (n_545, a[4], n_486);
  nand eco42 (n_486, n_839, n_840);
  or eco43 (n_547, n_496, a[5]);
  or eco44 (n_549, b[7], wc10);
  or eco45 (n_535, wc8, a[6]);
  not eco46 (wc8, b[6]);
  or eco47 (n_534, b[6], wc9);
  not eco48 (wc9, a[6]);
  or eco49 (n_544, wc11, a[7]);
  not eco50 (wc10, a[7]);
  or eco51 (n_558, n_482, wc12);
  not eco52 (wc11, b[7]);
  nand eco53 (n_565, n_473, n_474);
  not eco54 (wc12, n_515);
  nand eco55 (n_569, n_489, n_490);
  nand eco56 (n_571, n_481, n_482);
  nand eco57 (n_573, n_505, n_506);
  or eco58 (n_803, patchNew_wc10, n_495);
  or eco59 (n_804, patchNew_n_451, wc17);
  nand eco60 (n_495, n_758, n_759);
  not eco61 (wc17, n_495);
  or eco62 (n_504, wc25, n_729);
  not eco63 (wc20, n_504);
  or eco64 (n_508, wc38, n_684);
  not eco65 (wc21, n_508);
  or eco66 (n_480, wc35, n_669);
  not eco67 (wc22, n_480);
  or eco68 (n_728, n_725, n_471);
  not eco69 (wc25, n_728);
  nand eco70 (n_729, n_726, n_727);
  or eco71 (n_488, wc29, n_714);
  nand eco72 (n_665, b[2], a[2]);
  or eco73 (n_837, wc52, b[3]);
  not eco74 (wc52, op[0]);
  or eco75 (n_840, op[0], wc55);
  or eco76 (n_838, op[0], wc53);
  or eco77 (n_726, wc28, op[1]);
  or eco78 (n_727, wc50, n_472);
  not eco79 (wc26, n_488);
  or eco80 (n_492, wc31, n_699);
  not eco81 (wc28, n_564);
  not eco82 (wc27, n_492);
  nand eco83 (n_564, n_827, n_828);
  or eco84 (n_713, n_710, n_471);
  not eco85 (wc29, n_713);
  nand eco86 (n_714, n_711, n_712);
  nand eco87 (n_572, n_829, n_830);
  nand eco88 (n_597, n_496, a[5]);
  nand eco89 (n_497, n_588, n_765);
  nand eco90 (n_827, n_503, n_497);
  nand eco91 (n_503, n_547, n_597);
  or eco92 (n_828, n_503, n_497);
  or eco93 (n_711, wc30, op[1]);
  or eco94 (n_712, wc48, n_472);
  or eco95 (n_517, n_636, n_516);
  or eco96 (n_636, n_635, wc32);
  nand eco97 (n_516, n_549, n_534);
  or eco98 (n_520, n_648, n_519);
  or eco99 (n_648, n_647, wc33);
  nand eco100 (n_519, n_544, n_535);
  not eco101 (wc30, n_572);
  or eco102 (n_698, n_695, n_471);
  not eco103 (wc31, n_698);
  nand eco104 (n_699, n_696, n_697);
  or eco105 (n_696, wc36, op[1]);
  nand eco106 (n_588, n_486, a[4]);
  nand eco107 (n_765, n_545, n_485);
  or eco108 (n_635, n_634, wc37);
  not eco109 (wc32, n_515);
  or eco110 (n_518, a[5], wc62);
  or eco111 (n_697, wc44, n_472);
  nand eco112 (n_485, n_591, n_768);
  or eco113 (n_647, n_646, wc34);
  not eco114 (wc33, n_518);
  not eco115 (wc35, n_668);
  nand eco116 (n_829, n_487, n_485);
  nand eco117 (n_487, n_545, n_588);
  or eco118 (n_830, n_487, n_485);
  nand eco119 (n_646, n_645, n_482);
  not eco120 (wc34, n_489);
  nand eco121 (n_570, n_831, n_832);
  nand eco122 (n_669, n_666, n_667);
  or eco123 (n_668, n_665, n_471);
  nand eco124 (n_591, n_483, a[3]);
  nand eco125 (n_768, n_542, n_484);
  not eco126 (wc36, n_570);
  nand eco127 (n_645, n_576, n_490);
  nand eco128 (n_634, n_633, n_481);
  not eco129 (wc37, n_490);
  or eco130 (n_683, n_680, n_471);
  not eco131 (wc38, n_683);
  nand eco132 (n_684, n_681, n_682);
  nand eco133 (n_633, n_575, n_489);
  or eco134 (n_666, wc39, op[1]);
  or eco135 (n_667, wc49, n_472);
  nand eco136 (n_585, n_475, a[2]);
  nand eco137 (n_484, n_585, n_762);
  nand eco138 (n_831, n_491, n_484);
  nand eco139 (n_491, n_542, n_591);
  or eco140 (n_832, n_491, n_484);
  nand eco141 (n_576, n_623, n_624);
  not eco142 (wc39, n_566);
  nand eco143 (n_762, n_541, n_479);
  or eco144 (n_681, wc40, op[1]);
  or eco145 (n_682, wc45, n_472);
  nand eco146 (n_575, n_614, n_615);
  nand eco147 (n_651, n_557, n_556);
  nand eco148 (n_566, n_833, n_834);
  nand eco149 (n_574, n_835, n_836);
  or eco150 (n_557, n_519, wc41);
  nand eco151 (n_556, n_516, n_544);
  not eco152 (wc40, n_574);
  not eco153 (wc41, n_603);
  nand eco154 (n_614, n_474, n_537);
  or eco155 (n_615, n_613, b[0]);
  nand eco156 (n_654, n_560, n_559);
  or eco157 (n_560, n_516, wc43);
  nand eco158 (n_559, n_519, n_549);
  nand eco159 (n_833, n_476, n_479);
  nand eco160 (n_476, n_541, n_585);
  nand eco161 (n_479, n_600, n_777);
  or eco162 (n_834, n_476, n_479);
  nand eco163 (n_623, n_473, n_539);
  or eco164 (n_624, n_622, wc42);
  nand eco165 (n_600, n_477, a[1]);
  nand eco166 (n_603, n_555, n_515);
  or eco167 (n_622, n_537, a[0]);
  not eco168 (wc42, b[0]);
  not eco169 (wc43, n_606);
  nand eco170 (n_777, n_478, n_543);
  nand eco171 (n_835, n_478, n_507);
  nand eco172 (n_478, n_581, n_582);
  nand eco173 (n_507, n_543, n_600);
  or eco174 (n_836, n_478, n_507);
  or eco175 (n_613, n_539, wc47);
  not eco176 (wc44, n_569);
  nand eco177 (n_606, n_558, n_518);
  not eco178 (wc45, n_573);
  nand eco179 (n_472, op[1], op[0]);
  not eco180 (wc47, a[0]);
  not eco181 (wc48, n_571);
  or eco182 (n_758, n_582, n_471);
  nand eco183 (n_759, n_562, n_471);
  or eco184 (n_555, n_481, wc51);
  not eco185 (wc49, n_565);
  nand eco186 (n_562, n_841, n_842);
  or eco187 (n_471, wc68, op[0]);
  nand eco188 (n_582, a[0], b[0]);
  nand eco189 (n_710, b[4], a[4]);
  not eco190 (wc50, n_563);
  nand eco191 (n_725, b[5], a[5]);
  nand eco192 (n_563, n_515, n_518);
  nand eco193 (n_680, b[1], a[1]);
  or eco194 (n_581, b[0], wc63);
  nand eco195 (n_695, b[3], a[3]);
  not eco196 (wc53, b[3]);
  not eco197 (wc51, n_518);
  or eco198 (n_839, wc54, b[4]);
  not eco199 (wc54, op[0]);
  not eco200 (wc55, b[4]);
  or eco201 (n_842, a[0], wc57);
  or eco202 (n_841, wc56, b[0]);
  not eco203 (wc56, a[0]);
  not eco204 (wc57, b[0]);
  or eco205 (n_846, op[0], wc61);
  or eco206 (n_845, wc60, b[5]);
  not eco207 (wc60, op[0]);
  not eco208 (wc61, b[5]);
  not eco209 (wc62, b[5]);
  or eco210 (n_849, wc64, b[1]);
  not eco211 (wc63, op[0]);
  or eco212 (n_850, op[0], wc65);
  not eco213 (wc64, op[0]);
  not eco214 (wc65, b[1]);
  not eco215 (wc68, op[1]);
  or eco216 (n_851, wc66, b[2]);
  not eco217 (wc66, op[0]);
  or eco218 (n_852, op[0], wc67);
  not eco219 (wc67, b[2]);
  not eco220 (wc69, n_651);
  not eco221 (wc70, n_654);
  or eco222 (patchNew_n_69, patchNew_n_505, patchNew_n_264);
  not eco223 (patchNew_wc66, patchNew_n_69);
  not eco224 (patchNew_wc63, patchNew_n_69);
  not eco225 (patchNew_wc68, patchNew_n_69);
  not eco226 (patchNew_wc67, patchNew_n_69);
  not eco227 (patchNew_wc65, patchNew_n_69);
  not eco228 (patchNew_wc69, patchNew_n_69);
  not eco229 (patchNew_wc10, patchNew_n_451);
  nand eco230 (patchNew_n_451, patchNew_n_804, patchNew_n_805);
  or eco231 (patchNew_n_804, patchNew_wc12, patchNew_n_450);
  or eco232 (patchNew_n_805, patchNew_n_502, patchNew_wc13);
  nand eco233 (patchNew_n_505, patchNew_n_455, patchNew_n_705);
  or eco234 (patchNew_n_264, wc52, op[1]);
  not eco235 (patchNew_wc12, patchNew_n_502);
  nand eco236 (patchNew_n_450, patchNew_n_811, patchNew_n_812);
  nand eco237 (patchNew_n_502, patchNew_n_806, patchNew_n_807);
  not eco238 (patchNew_wc13, patchNew_n_450);
  or eco239 (patchNew_n_806, wc20, n_480);
  or eco240 (patchNew_n_807, n_504, wc22);
  or eco241 (patchNew_n_811, patchNew_wc17, n_488);
  or eco242 (patchNew_n_812, patchNew_n_503, wc26);
  not eco243 (patchNew_wc17, patchNew_n_503);
  nand eco244 (patchNew_n_503, patchNew_n_819, patchNew_n_820);
  or eco245 (patchNew_n_819, wc27, n_508);
  or eco246 (patchNew_n_820, n_492, wc21);
  or eco247 (patchNew_n_455, wc7, b[5]);
  nand eco248 (patchNew_n_705, patchNew_n_475, patchNew_n_413);
  or eco249 (patchNew_n_475, wc61, a[5]);
  nand eco250 (patchNew_n_413, patchNew_n_522, patchNew_n_687);
  or eco251 (patchNew_n_522, wc3, b[4]);
  nand eco252 (patchNew_n_687, n_482, patchNew_n_369);
  nand eco253 (patchNew_n_369, n_490, patchNew_n_657);
  nand eco254 (patchNew_n_657, n_489, patchNew_n_410);
  nand eco255 (patchNew_n_410, patchNew_n_521, patchNew_n_615);
  or eco256 (patchNew_n_521, wc1, b[2]);
  nand eco257 (patchNew_n_615, n_474, patchNew_n_360);
  nand eco258 (patchNew_n_360, n_506, patchNew_n_579);
  nand eco259 (patchNew_n_579, n_505, patchNew_n_496);
  or eco260 (patchNew_n_496, wc42, a[0]);
endmodule