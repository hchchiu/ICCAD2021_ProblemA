module top(o, a, b, c);
output o;
input a, b, c;
AND g1(o, a, b, c);
endmodule
