module top_eco(n_594, clk,\op[0] ,\a[0] ,\a[1] ,\a[5] ,\b[0] ,\b[1] ,\b[2] ,\b[3] ,\b[5] ,\op[1] , n_523, n_568, wc1, n_522, n_525, n_534, n_569, n_570, wc8, n_571, n_590, n_596, n_545, n_558, n_521, n_554, n_739, n_718, n_551, n_593, n_676, n_539, n_780, wc52, wc54, wc55, wc56, wc58, parity, overflow, greater,\y[0] , is_eq,\y[1] ,\y[2] ,\y[3] ,\y[4] ,\y[5] ,\y[6] ,\y[7] , less);
  input n_594, clk,\op[0] ,\a[0] ;
  input \a[1] ,\a[5] ,\b[0] ,\b[1] ,\b[2] ;
  input \b[3] ,\b[5] ,\op[1] , n_523, n_568;
  input wc1, n_522, n_525, n_534, n_569;
  input n_570, wc8, n_571, n_590, n_596;
  input n_545, n_558, n_521, n_554, n_739;
  input n_718, n_551, n_593, n_676, n_539;
  input n_780, wc52, wc54, wc55, wc56;
  input wc58;
  output parity, overflow, greater,\y[0] ;
  output is_eq,\y[1] ,\y[2] ,\y[3] ,\y[4] ;
  output \y[5] ,\y[6] ,\y[7] , less;
  wire nadd_28_29_n_21, nwc7, nn_503, nn_113;
  wire nn_292, nlt_44_17_n_37, nn_295, nwc0, nn_121;
  wire nn_296, nn_298, nn_301, nsub_33_29_n_54, nlt_44_17_n_71;
  wire nn_276, nn_505, nwc3, nn_110, nn_241;
  wire nn_504, nwc4, nn_506, nwc5, ntemp_y5;
  wire ntemp_y0, nn_495, nwc6, nn_510, nn_496;
  wire nn_508, nn_426, ngt_43_12_n_36, nn_258, nn_109;
  wire nn_242, nn_509, nwc8, ntemp_y4, nwc9;
  wire ntemp_y1, nn_489, nn_511, nwc10, nn_513;
  wire nwc11, ntemp_y2, ntemp_y3, nn_514, nwc12;
  wire nwc13, nn_283, nn_483, nn_484, nn_521;
  wire nn_490, nn_477, nn_478, nn_253, nwc14;
  wire nn_287, nwc15, nn_281, nwc16, nn_252;
  wire nn_456, nn_457, nn_472, nwc17, nn_278;
  wire nn_450, nsub_33_29_n_67, nn_522, nn_451, nn_524;
  wire nwc18, nadd_28_29_n_60, nn_525, nwc19, nn_462;
  wire nn_463, nn_358, nn_468, nn_469, nwc20;
  wire nn_254, nwc21, nn_257, nn_418, nlt_44_17_n_36;
  wire nlt_44_17_n_88, nn_442, nwc22, nn_427, nn_306;
  wire nn_360, nwc44, nn_361, nn_362, nn_438;
  wire nn_439, nn_445, nn_255, nwc23, nn_285;
  wire nn_318, nn_421, nlt_44_17_n_44, nn_294, nlt_44_17_n_87;
  wire nadd_28_29_n_47, nadd_28_29_n_50, nwc25, nn_289, nn_300;
  wire ngt_43_12_n_87, nn_527, nwc26, nadd_28_29_n_56, nn_528;
  wire nwc27, nn_432, nn_433, nn_529, nwc28;
  wire nn_530, nn_531, nn_532, nn_533, nsub_33_29_n_63;
  wire nn_534, nn_397, nn_244, nlt_44_17_n_66, nn_412;
  wire nn_402, nn_403, nn_394, ngt_43_12_n_66, nn_409;
  wire nn_406, nn_299, ngt_43_12_n_65, nn_293, nlt_44_17_n_65;
  wire nadd_28_29_n_41, nsub_33_29_n_48, nn_290, nn_260, nn_535;
  wire nn_536, nwc30, nn_259, nn_537, nwc31;
  wire nn_538, nwc32, nn_243, nn_539, nsub_33_29_n_32;
  wire nsub_33_29_n_60, nn_540, nn_541, nwc34, nadd_28_29_n_53;
  wire nn_542, nwc35, nn_325, nn_502, nn_363;
  wire nn_499, nn_369, nn_370, nn_381, nn_382;
  wire nn_390, nn_391, nn_375, nn_376, nn_280;
  wire nn_286, nwc36, nwc37, nn_359, nn_249;
  wire nn_284, ngt_43_12_n_34, nn_297, nn_288, nn_282;
  wire nn_389, nn_354, nn_355, nn_330, nn_331;
  wire nn_342, nn_343, nn_348, nn_349, nn_368;
  wire nwc39, nn_543, nwc40, nn_544, nwc41;
  wire nwc43, nwc42, nn_364, nn_336, nn_337;
  wire nwc55, nwc45, nadd_28_29_n_51, nwc46, nn_312;
  wire nn_310, nlt_44_17_n_68, nwc51, nwc52, nwc53;
  wire nwc54, nwc56, nwc57, nn_346, nn_347;
  wire nn_34, nn_308, nn_307, nn_27, nn_24;
  wire nadd_28_29_n_45, nn_323, nn_317, nn_320, nwc58;
  wire nn_332, nn_262, nadd_28_29_n_44, nwc65, nwc66;
  wire nn_415, nwc67;
  nand eco1 (nadd_28_29_n_21,\a[0] , nn_113);
  nand eco2 (parity, nn_503, nn_504);
  assign overflow = \y[7] ;
  not eco4 (greater, ngt_43_12_n_36);
  and eco5 (\y[0] , ntemp_y0, nwc53);
  and eco6 (is_eq, ngt_43_12_n_36, nlt_44_17_n_36);
  and eco7 (\y[1] , ntemp_y1, nwc52);
  and eco8 (\y[2] , nwc54, ntemp_y2);
  and eco9 (\y[3] , nwc55, ntemp_y3);
  and eco10 (\y[4] , nwc56, ntemp_y4);
  and eco11 (\y[5] , nwc57, ntemp_y5);
  nor eco12 (\y[6] , nn_472, nn_358);
  not eco13 (\y[7] , nn_358);
  and eco14 (less, ngt_43_12_n_36, nwc51);
  not eco15 (nwc7, nn_242);
  or eco16 (nn_503, nwc3, nn_110);
  nand eco17 (nn_113, nn_306, nn_360);
  nand eco18 (nn_292, nn_113, nlt_44_17_n_37);
  not eco19 (nlt_44_17_n_37,\a[0] );
  or eco20 (nn_295, nwc0,\a[1] );
  not eco21 (nwc0, nn_121);
  nand eco22 (nn_121, nn_361, nn_362);
  or eco23 (nn_296, nn_121,\a[1] );
  or eco24 (nn_298, nn_113, wc52);
  nand eco25 (nn_301, nsub_33_29_n_54, nlt_44_17_n_71);
  nand eco26 (nsub_33_29_n_54, nlt_44_17_n_66, nn_412);
  not eco27 (nlt_44_17_n_71, nn_262);
  or eco28 (nn_276,\b[5] , wc58);
  or eco29 (nn_505, nwc5, ntemp_y5);
  not eco30 (nwc3, nn_241);
  nand eco31 (nn_110, nn_508, nn_509);
  nand eco32 (nn_241, nn_505, nn_506);
  or eco33 (nn_504, nn_241, nwc4);
  not eco34 (nwc4, nn_110);
  or eco35 (nn_506, ntemp_y0, nwc6);
  not eco36 (nwc5, ntemp_y0);
  nand eco37 (ntemp_y5, nn_495, nn_496);
  nand eco38 (ntemp_y0, nn_390, nn_391);
  or eco39 (nn_495,\op[1] , nwc13);
  not eco40 (nwc6, ntemp_y5);
  or eco41 (nn_510, nwc9, ntemp_y1);
  nand eco42 (nn_496, nn_284,\op[1] );
  or eco43 (nn_508, nwc7, nn_109);
  nand eco44 (nn_426, nadd_28_29_n_47, nadd_28_29_n_50);
  nand eco45 (ngt_43_12_n_36, n_593, nn_445);
  nand eco46 (nn_258, nn_533, nn_534);
  nand eco47 (nn_109, nn_513, nn_514);
  nand eco48 (nn_242, nn_510, nn_511);
  or eco49 (nn_509, nn_242, nwc8);
  not eco50 (nwc8, nn_109);
  nand eco51 (ntemp_y4, nn_489, nn_490);
  not eco52 (nwc9, ntemp_y4);
  nand eco53 (ntemp_y1, nn_438, nn_439);
  or eco54 (nn_489,\op[1] , nwc14);
  or eco55 (nn_511, ntemp_y4, nwc10);
  not eco56 (nwc10, ntemp_y1);
  or eco57 (nn_513, nwc11, ntemp_y2);
  not eco58 (nwc11, ntemp_y3);
  nand eco59 (ntemp_y2, nn_462, nn_463);
  nand eco60 (ntemp_y3, nn_483, nn_484);
  or eco61 (nn_514, ntemp_y3, nwc12);
  not eco62 (nwc12, ntemp_y2);
  not eco63 (nwc13, nn_283);
  nand eco64 (nn_283, nn_477, nn_478);
  or eco65 (nn_483,\op[1] , nwc15);
  nand eco66 (nn_484, nn_282,\op[1] );
  nand eco67 (nn_521, nsub_33_29_n_67, n_558);
  nand eco68 (nn_490, nn_288,\op[1] );
  or eco69 (nn_477, nwc16,\op[0] );
  nand eco70 (nn_478, nn_253,\op[0] );
  nand eco71 (nn_253, nn_521, nn_522);
  not eco72 (nwc14, nn_287);
  nand eco73 (nn_287, nn_456, nn_457);
  not eco74 (nwc15, nn_281);
  nand eco75 (nn_281, nn_450, nn_451);
  not eco76 (nwc16, nn_252);
  nand eco77 (nn_252, nn_524, nn_525);
  or eco78 (nn_456, nwc20,\op[0] );
  nand eco79 (nn_457, nn_255,\op[0] );
  or eco80 (nn_472, nwc17,\op[1] );
  not eco81 (nwc17, nn_278);
  or eco82 (nn_278, nwc22, nn_427);
  or eco83 (nn_450, nwc21,\op[0] );
  nand eco84 (nsub_33_29_n_67, n_521, nn_418);
  or eco85 (nn_522, nsub_33_29_n_67, n_558);
  nand eco86 (nn_451, nn_258,\op[0] );
  or eco87 (nn_524, nwc18, n_558);
  not eco88 (nwc18, nadd_28_29_n_60);
  nand eco89 (nadd_28_29_n_60, n_739, nn_421);
  or eco90 (nn_525, nadd_28_29_n_60, nwc19);
  not eco91 (nwc19, n_558);
  or eco92 (nn_462,\op[1] , nwc23);
  nand eco93 (nn_463, nn_286,\op[1] );
  or eco94 (nn_358, nn_468, nn_469);
  or eco95 (nn_468, nwc65,\op[1] );
  nand eco96 (nn_469,\op[0] , nlt_44_17_n_68);
  not eco97 (nwc20, nn_254);
  nand eco98 (nn_254, nn_529, nn_530);
  not eco99 (nwc21, nn_257);
  nand eco100 (nn_257, nn_527, nn_528);
  nand eco101 (nn_418, nsub_33_29_n_54, n_522);
  nand eco102 (nlt_44_17_n_36, nlt_44_17_n_88, nn_442);
  nand eco103 (nlt_44_17_n_88, nn_346, nn_347);
  nand eco104 (nn_442, nn_294, nlt_44_17_n_87);
  not eco105 (nwc22, nn_426);
  or eco106 (nn_427, nwc45,\op[0] );
  or eco107 (nn_306, wc8, clk);
  nand eco108 (nn_360,\b[0] , clk);
  not eco109 (nwc44,\a[0] );
  or eco110 (nn_361, wc1, clk);
  nand eco111 (nn_362,\b[1] , clk);
  or eco112 (nn_438,\op[1] , nwc25);
  nand eco113 (nn_439, nn_290,\op[1] );
  nand eco114 (nn_445, nn_300, ngt_43_12_n_87);
  nand eco115 (nn_255, nn_531, nn_532);
  not eco116 (nwc23, nn_285);
  nand eco117 (nn_285, nn_432, nn_433);
  or eco118 (nn_318, nn_121, wc54);
  nand eco119 (nn_421, nadd_28_29_n_47, n_590);
  or eco120 (nlt_44_17_n_44, wc55,\b[2] );
  nand eco121 (nn_294, nlt_44_17_n_66, nn_406);
  nor eco122 (nlt_44_17_n_87, nn_262, nn_307);
  nand eco123 (nadd_28_29_n_47, nadd_28_29_n_45, nn_415);
  and eco124 (nadd_28_29_n_50, nn_312, n_590);
  not eco125 (nwc25, nn_289);
  nand eco126 (nn_289, nn_402, nn_403);
  nand eco127 (nn_300, ngt_43_12_n_66, nn_409);
  nor eco128 (ngt_43_12_n_87, nn_332, nn_308);
  or eco129 (nn_527, nwc26, n_554);
  not eco130 (nwc26, nadd_28_29_n_56);
  nand eco131 (nadd_28_29_n_56, n_676, nn_397);
  or eco132 (nn_528, nadd_28_29_n_56, nwc27);
  not eco133 (nwc27, n_554);
  or eco134 (nn_432, nwc67,\op[0] );
  nand eco135 (nn_433, nn_244,\op[0] );
  or eco136 (nn_529, nwc28, n_545);
  not eco137 (nwc28, nadd_28_29_n_47);
  or eco138 (nn_530, nadd_28_29_n_47, nwc66);
  nand eco139 (nn_531, nsub_33_29_n_54, n_545);
  or eco140 (nn_532, nsub_33_29_n_54, n_545);
  nand eco141 (nn_533, nsub_33_29_n_63, n_554);
  nand eco142 (nsub_33_29_n_63, nlt_44_17_n_44, nn_394);
  or eco143 (nn_534, nsub_33_29_n_63, n_554);
  nand eco144 (nn_397, nadd_28_29_n_41, n_596);
  nand eco145 (nn_244, nn_535, nn_536);
  nand eco146 (nlt_44_17_n_66, nn_24, n_523);
  nand eco147 (nn_412, nsub_33_29_n_48, nlt_44_17_n_65);
  or eco148 (nn_402, nwc30,\op[0] );
  nand eco149 (nn_403, nn_260,\op[0] );
  nand eco150 (nn_394, nsub_33_29_n_48, n_525);
  nand eco151 (ngt_43_12_n_66, nn_27, nn_310);
  nand eco152 (nn_409, nn_299, ngt_43_12_n_65);
  nand eco153 (nn_406, nn_293, nlt_44_17_n_65);
  nand eco154 (nn_299, nn_381, nn_382);
  not eco155 (ngt_43_12_n_65, nn_24);
  nand eco156 (nn_293, nn_375, nn_376);
  not eco157 (nlt_44_17_n_65, nn_27);
  nand eco158 (nadd_28_29_n_41, nn_325, nn_502);
  nand eco159 (nsub_33_29_n_48, nn_318, nn_499);
  nand eco160 (nn_290, nn_369, nn_370);
  nand eco161 (nn_260, nn_539, nn_540);
  nand eco162 (nn_535, nsub_33_29_n_48, n_551);
  or eco163 (nn_536, nsub_33_29_n_48, n_551);
  not eco164 (nwc30, nn_259);
  nand eco165 (nn_259, nn_541, nn_542);
  or eco166 (nn_537, nwc31, n_551);
  not eco167 (nwc31, nadd_28_29_n_41);
  or eco168 (nn_538, nadd_28_29_n_41, nwc32);
  not eco169 (nwc32, n_551);
  nand eco170 (nn_243, nn_537, nn_538);
  nand eco171 (nn_539, nsub_33_29_n_32, nsub_33_29_n_60);
  nand eco172 (nsub_33_29_n_32, nlt_44_17_n_37, nn_113);
  nand eco173 (nsub_33_29_n_60, nn_318, nn_295);
  or eco174 (nn_540, nsub_33_29_n_32, nsub_33_29_n_60);
  or eco175 (nn_541, nwc34, nadd_28_29_n_53);
  not eco176 (nwc34, nadd_28_29_n_21);
  nand eco177 (nadd_28_29_n_53, nn_296, nn_325);
  or eco178 (nn_542, nadd_28_29_n_21, nwc35);
  not eco179 (nwc35, nadd_28_29_n_53);
  nand eco180 (nn_325, nn_121,\a[1] );
  or eco181 (nn_502, nwc36, nadd_28_29_n_21);
  or eco182 (nn_363,\a[1] ,\a[0] );
  nand eco183 (nn_499, nn_295, nsub_33_29_n_32);
  or eco184 (nn_369, nn_368, nwc39);
  nand eco185 (nn_370, nn_249,\op[0] );
  nand eco186 (nn_381, nn_298, ngt_43_12_n_34);
  nand eco187 (nn_382, nn_297, nn_121);
  or eco188 (nn_390, nn_389, nn_113);
  nand eco189 (nn_391, nn_280, nn_113);
  nand eco190 (nn_375, nn_292,\a[1] );
  or eco191 (nn_376, nwc37, nn_121);
  nand eco192 (nn_280, nn_330, nn_331);
  nand eco193 (nn_286, nn_348, nn_349);
  not eco194 (nwc36, nn_296);
  not eco195 (nwc37, nn_359);
  or eco196 (nn_359, nn_363, nwc42);
  nand eco197 (nn_249, nn_543, nn_544);
  nand eco198 (nn_284, nn_342, nn_343);
  not eco199 (ngt_43_12_n_34,\a[1] );
  or eco200 (nn_297, nn_364, nn_113);
  nand eco201 (nn_288, nn_354, nn_355);
  nand eco202 (nn_282, nn_336, nn_337);
  nand eco203 (nn_389,\a[0] , n_539);
  or eco204 (nn_354,\op[0] , n_739);
  nand eco205 (nn_355, n_545,\op[0] );
  or eco206 (nn_330, n_539, nwc44);
  or eco207 (nn_331, nwc43,\a[0] );
  or eco208 (nn_342,\op[0] , n_780);
  nand eco209 (nn_343, n_558,\op[0] );
  or eco210 (nn_348,\op[0] , n_676);
  nand eco211 (nn_349, n_551,\op[0] );
  or eco212 (nn_368, nwc46,\op[0] );
  not eco213 (nwc39, nn_121);
  or eco214 (nn_543, nwc40, nn_121);
  not eco215 (nwc40,\a[1] );
  or eco216 (nn_544,\a[1] , nwc41);
  not eco217 (nwc41, nn_121);
  not eco218 (nwc43, n_539);
  not eco219 (nwc42, nn_113);
  nand eco220 (nn_364,\a[1] ,\a[0] );
  or eco221 (nn_336,\op[0] , n_718);
  nand eco222 (nn_337, n_554,\op[0] );
  not eco223 (nwc55, nn_358);
  not eco224 (nwc45, nadd_28_29_n_51);
  nand eco225 (nadd_28_29_n_51, nn_312, nn_320);
  not eco226 (nwc46,\a[1] );
  or eco227 (nn_312,\b[5] ,\a[5] );
  or eco228 (nn_310,\b[3] , wc56);
  not eco229 (nlt_44_17_n_68, nn_34);
  not eco230 (nwc51, nlt_44_17_n_36);
  not eco231 (nwc52, nn_358);
  not eco232 (nwc53, nn_358);
  not eco233 (nwc54, nn_358);
  not eco234 (nwc56, nn_358);
  not eco235 (nwc57, nn_358);
  or eco236 (nn_346, nn_34, nn_308);
  nand eco237 (nn_347, n_569, nn_307);
  nand eco238 (nn_34, nn_317, nn_276);
  nand eco239 (nn_308, n_569, n_571);
  nand eco240 (nn_307, n_568, n_570);
  nand eco241 (nn_27, n_523, n_525);
  nand eco242 (nn_24, nn_310, nlt_44_17_n_44);
  nand eco243 (nadd_28_29_n_45, n_594, nn_323);
  nand eco244 (nn_323, n_676, n_718);
  or eco245 (nn_317, n_521, nwc58);
  nand eco246 (nn_320, n_739, n_780);
  not eco247 (nwc58, n_534);
  nand eco248 (nn_332, n_521, nn_276);
  nand eco249 (nn_262, n_522, n_534);
  and eco250 (nadd_28_29_n_44, n_594, n_596);
  not eco251 (nwc65, nn_301);
  not eco252 (nwc66, n_545);
  nand eco253 (nn_415, nadd_28_29_n_41, nadd_28_29_n_44);
  not eco254 (nwc67, nn_243);
endmodule
