module top_eco(n17, n25, n145, n146, n148, n124, n125, n127, n130, n131, n133, n136, n137, n138, n142, n144, n407, n155, n157, n161, n164, n165, n168, n174, n179, n195, n197, n200, n204, n207, n211, n261, n262, n264, n330, n331, n332, n334, n342, n374, n375, n376, n378, n389, n397, n921, n928, n439, n444, n473, n476, n477, n478, n479, n487, n496, n511, n512, n514, n515, n530, n533, n535, n540, n541, n547, n557, n586, n587, n589, n613, n624, n625, n630, n634, n638, n642, n660, n661, n663, n666, n667, n669, n673, n674, n676, n677, n679, n682, n683, n685, n692, n694, n698, n701, n702, n705, n711, n712, n713, n717, n721, n727, n732, n735, n739, n742, n756, n761, n762, n774, n781, n782, n785, n790, n793, n804, n822, n834, n846, n854, n858, n864, n866, n867, n887, n890, n891, n894, n906, n909, n1962, n935, n941, n951, n952, n953, n1004, n1011, n1012, n1053, n1056, n1059, n1066, n1070, n1075, n1076, n1094, n1095, n1106, n1112, n1113, n1115, n1126, n1131, n1147, n1154, n1168, n1193, n1204, n1206, n1255, n1308, n1336, n1375, n1381, n1386, n1407, n1423, n1424, n1453, n1454, n1461, n1515, n1530, n1546, n1555, n1562, n1574, n1597, n1614, n1627, n1666, n1699, n1702, n1708, n1710, n1717, n1718, n1723, n1754, n1778, n1897, n2007, g48, n69, n74, n75, n76, n84, n2015, n1808, n1819, n1833, n1844, n1851, n1866, n1891, n1910, n1921, n1949, n1955, n1972, n1960, n1965, n1967, n1602, n1604, n1620, n1622, n1824, n1826, n1835, n1837, n1856, n1859, n1873, n1875, n1933, n1940, n1942);
  input n17, n25, n145, n146;
  input n148, n124, n125, n127, n130;
  input n131, n133, n136, n137, n138;
  input n142, n144, n407, n155, n157;
  input n161, n164, n165, n168, n174;
  input n179, n195, n197, n200, n204;
  input n207, n211, n261, n262, n264;
  input n330, n331, n332, n334, n342;
  input n374, n375, n376, n378, n389;
  input n397, n921, n928, n439, n444;
  input n473, n476, n477, n478, n479;
  input n487, n496, n511, n512, n514;
  input n515, n530, n533, n535, n540;
  input n541, n547, n557, n586, n587;
  input n589, n613, n624, n625, n630;
  input n634, n638, n642, n660, n661;
  input n663, n666, n667, n669, n673;
  input n674, n676, n677, n679, n682;
  input n683, n685, n692, n694, n698;
  input n701, n702, n705, n711, n712;
  input n713, n717, n721, n727, n732;
  input n735, n739, n742, n756, n761;
  input n762, n774, n781, n782, n785;
  input n790, n793, n804, n822, n834;
  input n846, n854, n858, n864, n866;
  input n867, n887, n890, n891, n894;
  input n906, n909, n1962, n935, n941;
  input n951, n952, n953, n1004, n1011;
  input n1012, n1053, n1056, n1059, n1066;
  input n1070, n1075, n1076, n1094, n1095;
  input n1106, n1112, n1113, n1115, n1126;
  input n1131, n1147, n1154, n1168, n1193;
  input n1204, n1206, n1255, n1308, n1336;
  input n1375, n1381, n1386, n1407, n1423;
  input n1424, n1453, n1454, n1461, n1515;
  input n1530, n1546, n1555, n1562, n1574;
  input n1597, n1614, n1627, n1666, n1699;
  input n1702, n1708, n1710, n1717, n1718;
  input n1723, n1754, n1778, n1897, n2007;
  output g48, n69, n74, n75;
  output n76, n84, n2015, n1808, n1819;
  output n1833, n1844, n1851, n1866, n1891;
  output n1910, n1921, n1949, n1955, n1972;
  output n1960, n1965, n1967, n1602, n1604;
  output n1620, n1622, n1824, n1826, n1835;
  output n1837, n1856, n1859, n1873, n1875;
  output n1933, n1940, n1942;
  buf eco1 (n69, patchNew_n1959);
  buf eco2 (n74, patchNew_n2005);
  buf eco3 (n75, patchNew__xnor_GATE_0);
  buf eco4 (n76, patchNew_n2043);
  buf eco5 (n84, patchNew_n1913);
  nor eco6 (n2015, patchNew_n1945, patchNew_n1946);
  nor eco7 (n1808, patchNew_n1948, patchNew_n1949);
  nor eco8 (n1819, patchNew_n1964_n1886_29, patchNew__xnor_GATE_3);
  nor eco9 (n1833, patchNew_n1969, patchNew_n1063);
  nor eco10 (n1844, patchNew_n1983, patchNew_n1911);
  nor eco11 (n1851, patchNew_n1988, patchNew_n1989);
  nor eco12 (n1866, patchNew_n1994, patchNew_n1997);
  nor eco13 (n1891, patchNew_n2026, patchNew_n2028);
  nor eco14 (n1910, patchNew_n2046, patchNew_n2050);
  nor eco15 (n1921, patchNew_n2066_n2067_30, patchNew__xor_GATE_1);
  nor eco16 (n1949, patchNew_n2071_n2072_31, patchNew_n844);
  nor eco17 (n1955, patchNew_n2082, n1702);
  nor eco18 (n1972, patchNew_n2099, patchNew_n1791);
  and eco19 (n1824, patchNew_n1923, patchNew__xnor_GATE_2);
  and eco20 (n1826, patchNew_n1926, patchNew_n1860);
  and eco21 (n1856, patchNew_n1937, patchNew_n1907);
  and eco22 (n1859, patchNew_n1939, patchNew_n1940);
  and eco23 (n1602, patchNew_n1077, patchNew_n1717);
  and eco24 (n1604, patchNew_n1719, patchNew_n1720);
  and eco25 (n1835, patchNew_n1936, patchNew_n1976);
  and eco26 (n1837, patchNew_n1978, patchNew_n1979);
  and eco27 (n1873, patchNew_n1931, patchNew_n2010);
  and eco28 (n1875, patchNew_n2012, patchNew_n2009);
  not eco29 (n1933, patchNew__xnor_GATE_4);
  not eco30 (n1940, patchNew_n2058);
  or eco31 (n1942, patchNew_n2058, patchNew__xnor_GATE_4);
  not eco32 (n1960, patchNew__xnor_GATE_5);
  not eco33 (n1965, patchNew_n848);
  or eco34 (n1967, patchNew_n848, patchNew__xnor_GATE_5);
  and eco35 (n1620, patchNew_n1971, patchNew__xnor_GATE_6);
  and eco36 (n1622, patchNew_n2125, patchNew_n1972);
  buf eco37 (g48, 1'b0);
  or eco38 (patchNew_n1959, patchNew_new_n498_, patchNew_new_n499_);
  or eco39 (patchNew_n2005, patchNew_new_n514_, patchNew_new_n515_);
  nor eco40 (patchNew_n2043, patchNew_new_n536_, patchNew_new_n537_);
  or eco41 (patchNew_n1913, patchNew_new_n626_, patchNew_new_n629_);
  nor eco42 (patchNew_n844, patchNew_new_n255_, patchNew_new_n310_);
  nor eco43 (patchNew_n848, patchNew_new_n312_, patchNew_new_n313_);
  nor eco44 (patchNew_n1923, patchNew_new_n346_, patchNew_new_n631_);
  not eco45 (patchNew_n1926, patchNew_n1923);
  and eco46 (patchNew_n1931, patchNew__not_GATE_47, patchNew_new_n335_);
  not eco47 (patchNew_n1936, patchNew_n1978);
  not eco48 (patchNew_n1937, patchNew_n1939);
  nor eco49 (patchNew_n1939, patchNew_n1978, patchNew_new_n633_);
  not eco50 (patchNew_n1940, patchNew_n1907);
  and eco51 (patchNew_n1945, patchNew__not_GATE_156, patchNew_new_n638_);
  or eco52 (patchNew_n1946, patchNew_new_n640_, patchNew_new_n641_);
  nor eco53 (patchNew_n1948, patchNew_new_n635_, patchNew_new_n643_);
  nor eco54 (patchNew_n1949, patchNew_new_n274_, patchNew_new_n275_);
  or eco55 (patchNew_n1063, patchNew_new_n339_, patchNew_new_n340_);
  not eco56 (patchNew_n1077, patchNew_n1719);
  not eco57 (patchNew_n1717, patchNew_n1720);
  nor eco58 (patchNew_n1719, patchNew_n1946, patchNew_new_n646_);
  and eco59 (patchNew_n1720, n1255, patchNew__not_GATE_154);
  or eco60 (patchNew_n1791, patchNew__not_GATE_133, patchNew_new_n572_);
  not eco61 (patchNew_n1860, patchNew__xnor_GATE_2);
  nor eco62 (patchNew_n1907, patchNew_new_n544_, patchNew_new_n612_);
  and eco63 (patchNew_n1911, patchNew_new_n611_, patchNew__not_GATE_152);
  nor eco64 (patchNew_n1964_n1886_29, patchNew_new_n614_, patchNew_new_n649_);
  or eco65 (patchNew_n1969, patchNew_new_n648_, patchNew_new_n651_);
  not eco66 (patchNew_n1971, patchNew_n1972);
  and eco67 (patchNew_n1972, patchNew_n1949, patchNew_new_n346_);
  not eco68 (patchNew_n1976, patchNew_n1979);
  and eco69 (patchNew_n1978, patchNew__not_GATE_48, patchNew_new_n337_);
  nor eco70 (patchNew_n1979, patchNew_new_n653_, patchNew_new_n654_);
  or eco71 (patchNew_n1983, patchNew__not_GATE_160, patchNew_new_n656_);
  or eco72 (patchNew_n1988, patchNew_new_n611_, patchNew_new_n658_);
  nor eco73 (patchNew_n1989, patchNew_new_n287_, patchNew_new_n288_);
  and eco74 (patchNew_n1994, patchNew_new_n610_, patchNew__not_GATE_161);
  or eco75 (patchNew_n1997, patchNew_new_n301_, patchNew_new_n662_);
  not eco76 (patchNew_n2009, patchNew_n2010);
  nor eco77 (patchNew_n2010, patchNew_new_n664_, patchNew_new_n665_);
  not eco78 (patchNew_n2012, patchNew_n1931);
  nor eco79 (patchNew_n2026, patchNew_new_n608_, patchNew_new_n667_);
  or eco80 (patchNew_n2028, patchNew__not_GATE_163, patchNew_new_n605_);
  and eco81 (patchNew_n2046, patchNew_new_n602_, patchNew__not_GATE_164);
  or eco82 (patchNew_n2050, patchNew_new_n323_, patchNew_new_n598_);
  or eco83 (patchNew_n2058, patchNew_new_n308_, patchNew_new_n309_);
  nor eco84 (patchNew_n2066_n2067_30, patchNew_new_n594_, patchNew_new_n678_);
  nor eco85 (patchNew_n2071_n2072_31, patchNew_new_n681_, patchNew_new_n682_);
  or eco86 (patchNew_n2082, patchNew_new_n577_, patchNew_new_n688_);
  nor eco87 (patchNew_n2099, n1723, patchNew_new_n690_);
  not eco88 (patchNew_n2125, patchNew__xnor_GATE_6);
  not eco89 (patchNew__not_GATE_40, n1555);
  not eco90 (patchNew__not_GATE_81, patchNew_new_n436_);
  not eco91 (patchNew__not_GATE_37, n1453);
  nor eco92 (patchNew_new_n301_, patchNew_new_n299_, patchNew_new_n300_);
  and eco93 (patchNew_new_n271_, n211, patchNew__not_GATE_22);
  and eco94 (patchNew_new_n381_, n864, patchNew__not_GATE_62);
  not eco95 (patchNew__not_GATE_33, patchNew_new_n294_);
  not eco96 (patchNew__not_GATE_8, n541);
  nor eco97 (patchNew_new_n320_, n1546, patchNew_new_n319_);
  nor eco98 (patchNew_new_n382_, n867, n864);
  nor eco99 (patchNew_new_n242_, patchNew_new_n239_, patchNew_new_n241_);
  and eco100 (patchNew_new_n378_, n822, patchNew__not_GATE_60);
  and eco101 (patchNew_new_n434_, patchNew_new_n388_, patchNew_new_n433_);
  not eco102 (patchNew__not_GATE_21, patchNew_new_n269_);
  nor eco103 (patchNew_new_n309_, n1407, patchNew__xor_GATE_1);
  not eco104 (patchNew__not_GATE_39, n1423);
  and eco105 (patchNew_new_n262_, patchNew_new_n246_, patchNew__not_GATE_15);
  nor eco106 (patchNew_new_n335_, patchNew_new_n330_, patchNew_new_n334_);
  not eco107 (patchNew__not_GATE_22, patchNew_new_n270_);
  and eco108 (patchNew_new_n250_, patchNew__not_GATE_10, n547);
  nor eco109 (patchNew_new_n387_, patchNew_new_n380_, patchNew_new_n381_);
  not eco110 (patchNew__not_GATE_32, patchNew_new_n293_);
  nor eco111 (patchNew_new_n263_, patchNew_new_n244_, patchNew_new_n262_);
  and eco112 (patchNew_new_n321_, patchNew__not_GATE_40, patchNew_new_n319_);
  nor eco113 (patchNew_new_n484_, patchNew_new_n437_, patchNew_new_n483_);
  nor eco114 (patchNew_new_n362_, patchNew_new_n350_, patchNew_new_n361_);
  nor eco115 (patchNew_new_n350_, n739, n742);
  nor eco116 (patchNew_new_n383_, n781, n866);
  nor eco117 (patchNew_new_n334_, patchNew_new_n298_, patchNew_new_n301_);
  nor eco118 (patchNew_new_n273_, patchNew_new_n271_, patchNew_new_n272_);
  and eco119 (patchNew_new_n292_, patchNew__not_GATE_31, patchNew_new_n291_);
  and eco120 (patchNew_new_n373_, n756, patchNew_new_n372_);
  not eco121 (patchNew__not_GATE_105, patchNew_new_n507_);
  not eco122 (patchNew__not_GATE_77, patchNew_new_n420_);
  and eco123 (patchNew_new_n439_, patchNew__not_GATE_82, patchNew_new_n438_);
  and eco124 (patchNew_new_n277_, n625, patchNew_new_n263_);
  nor eco125 (patchNew_new_n261_, patchNew_new_n256_, patchNew_new_n260_);
  nor eco126 (patchNew_new_n304_, patchNew_new_n256_, patchNew_new_n303_);
  not eco127 (patchNew__not_GATE_17, patchNew_new_n264_);
  nor eco128 (patchNew_new_n450_, patchNew_new_n448_, patchNew_new_n449_);
  and eco129 (patchNew_new_n315_, patchNew__not_GATE_39, patchNew_n848);
  not eco130 (patchNew__not_GATE_41, patchNew_new_n246_);
  and eco131 (patchNew_new_n264_, n512, patchNew__not_GATE_16);
  and eco132 (patchNew_new_n371_, patchNew__not_GATE_59, patchNew_new_n369_);
  nor eco133 (patchNew_new_n279_, patchNew_new_n277_, patchNew_new_n278_);
  and eco134 (patchNew_new_n359_, n739, patchNew__not_GATE_54);
  and eco135 (patchNew_new_n394_, n953, n921);
  nor eco136 (patchNew_new_n251_, patchNew_new_n249_, patchNew_new_n250_);
  not eco137 (patchNew__not_GATE_52, n721);
  nor eco138 (patchNew_new_n398_, patchNew_new_n396_, patchNew_new_n397_);
  and eco139 (patchNew_new_n280_, patchNew__not_GATE_25, patchNew_new_n279_);
  not eco140 (patchNew__not_GATE_15, patchNew_new_n261_);
  not eco141 (patchNew__not_GATE_97, patchNew_new_n485_);
  and eco142 (patchNew_new_n241_, n557, patchNew__not_GATE_6);
  and eco143 (patchNew_new_n291_, patchNew__not_GATE_30, n1530);
  not eco144 (patchNew__not_GATE_30, n1562);
  not eco145 (patchNew__not_GATE_79, n887);
  nor eco146 (patchNew_new_n360_, patchNew_new_n350_, patchNew_new_n359_);
  and eco147 (patchNew_new_n312_, n1515, patchNew__not_GATE_38);
  nor eco148 (patchNew_new_n443_, patchNew_new_n441_, patchNew_new_n442_);
  and eco149 (patchNew_new_n352_, n732, n735);
  and eco150 (patchNew_new_n386_, patchNew__not_GATE_63, patchNew_new_n385_);
  and eco151 (patchNew_new_n339_, patchNew__not_GATE_49, patchNew_new_n268_);
  and eco152 (patchNew_new_n249_, patchNew_n499, patchNew__not_GATE_9);
  and eco153 (patchNew_new_n275_, patchNew__not_GATE_24, patchNew_new_n273_);
  not eco154 (patchNew__not_GATE_13, patchNew_new_n242_);
  and eco155 (patchNew_new_n397_, n909, n906);
  and eco156 (patchNew_new_n441_, n951, patchNew__not_GATE_84);
  not eco157 (patchNew__not_GATE_61, n858);
  not eco158 (patchNew__not_GATE_86, n1112);
  nor eco159 (patchNew_new_n246_, patchNew_new_n244_, patchNew_new_n245_);
  not eco160 (patchNew__not_GATE_9, n547);
  nor eco161 (patchNew_new_n393_, patchNew_new_n391_, patchNew_new_n392_);
  nor eco162 (patchNew_new_n438_, patchNew_new_n423_, patchNew_new_n437_);
  nor eco163 (patchNew_new_n472_, patchNew_new_n454_, patchNew__xnor_GATE_9);
  nor eco164 (patchNew_new_n396_, n894, patchNew_new_n395_);
  and eco165 (patchNew_new_n459_, n1112, patchNew__not_GATE_89);
  and eco166 (patchNew_new_n337_, patchNew_n1989, patchNew_n1931);
  nor eco167 (patchNew_new_n406_, patchNew_new_n394_, patchNew_new_n405_);
  and eco168 (patchNew_new_n452_, patchNew__not_GATE_86, patchNew_new_n450_);
  and eco169 (patchNew_new_n294_, n1308, patchNew__not_GATE_32);
  and eco170 (patchNew_new_n284_, n332, patchNew__not_GATE_28);
  not eco171 (patchNew__not_GATE_96, patchNew_new_n446_);
  not eco172 (patchNew__not_GATE_12, n586);
  nor eco173 (patchNew_new_n296_, n1530, patchNew_new_n295_);
  and eco174 (patchNew_new_n243_, patchNew__not_GATE_7, patchNew_new_n242_);
  and eco175 (patchNew_new_n230_, n331, patchNew__not_GATE_0);
  nor eco176 (patchNew_new_n318_, patchNew_new_n309_, patchNew_new_n317_);
  nor eco177 (patchNew_new_n254_, patchNew_new_n252_, patchNew_new_n253_);
  not eco178 (patchNew__not_GATE_60, patchNew_n1390);
  and eco179 (patchNew_new_n380_, patchNew_n1224, patchNew__not_GATE_61);
  nor eco180 (patchNew_new_n504_, patchNew_new_n302_, patchNew_new_n334_);
  nor eco181 (patchNew_new_n385_, patchNew_new_n382_, patchNew_new_n383_);
  and eco182 (patchNew_new_n361_, patchNew__not_GATE_55, patchNew_new_n360_);
  nor eco183 (patchNew_new_n340_, n262, patchNew_new_n268_);
  nor eco184 (patchNew_new_n237_, patchNew_new_n234_, patchNew_new_n236_);
  nor eco185 (patchNew_new_n379_, n822, n804);
  and eco186 (patchNew_new_n421_, n951, patchNew__not_GATE_77);
  not eco187 (patchNew__not_GATE_47, patchNew_new_n333_);
  and eco188 (patchNew_new_n256_, patchNew__not_GATE_12, patchNew_new_n255_);
  and eco189 (patchNew_new_n252_, patchNew_new_n248_, patchNew_new_n251_);
  nor eco190 (patchNew_new_n248_, patchNew_new_n240_, patchNew_new_n247_);
  not eco191 (patchNew__not_GATE_6, patchNew_new_n240_);
  nor eco192 (patchNew_new_n433_, patchNew_new_n378_, patchNew_new_n432_);
  not eco193 (patchNew__not_GATE_38, patchNew_n844);
  and eco194 (patchNew_new_n364_, n713, patchNew_new_n362_);
  not eco195 (patchNew__not_GATE_48, patchNew_new_n286_);
  and eco196 (patchNew_new_n444_, patchNew_new_n418_, patchNew_new_n443_);
  nor eco197 (patchNew_new_n356_, patchNew_new_n354_, patchNew_new_n355_);
  not eco198 (patchNew__not_GATE_49, n261);
  not eco199 (patchNew__not_GATE_70, patchNew_new_n403_);
  and eco200 (patchNew_new_n272_, patchNew_n1008, patchNew_n989);
  and eco201 (patchNew_new_n384_, n781, n866);
  not eco202 (patchNew__not_GATE_20, n262);
  and eco203 (patchNew_new_n402_, n854, patchNew__not_GATE_68);
  nor eco204 (patchNew_new_n245_, n613, patchNew_new_n243_);
  not eco205 (patchNew__not_GATE_29, n375);
  nor eco206 (patchNew_new_n458_, patchNew_new_n456_, patchNew_new_n457_);
  and eco207 (patchNew_new_n447_, n1094, patchNew_new_n446_);
  nor eco208 (patchNew_new_n376_, n756, patchNew_new_n372_);
  and eco209 (patchNew_new_n432_, patchNew__not_GATE_80, patchNew_n1390);
  nor eco210 (patchNew_new_n399_, n953, patchNew_n1188);
  not eco211 (patchNew__not_GATE_31, patchNew_new_n290_);
  nor eco212 (patchNew_new_n299_, n444, patchNew_new_n279_);
  nor eco213 (patchNew_new_n298_, patchNew_new_n292_, patchNew_new_n297_);
  and eco214 (patchNew_new_n228_, patchNew_new_n226_, patchNew_new_n227_);
  and eco215 (patchNew_new_n281_, n630, patchNew__not_GATE_26);
  and eco216 (patchNew_new_n313_, n1962, patchNew_n844);
  and eco217 (patchNew_new_n342_, patchNew_n1978, patchNew_n1063);
  and eco218 (patchNew_new_n453_, n1113, patchNew__not_GATE_87);
  and eco219 (patchNew_new_n287_, patchNew__not_GATE_29, patchNew_new_n281_);
  not eco220 (patchNew__not_GATE_82, patchNew_new_n428_);
  and eco221 (patchNew_new_n255_, n1453, patchNew__not_GATE_11);
  nor eco222 (patchNew_new_n463_, patchNew_new_n461_, patchNew_new_n462_);
  not eco223 (patchNew__not_GATE_80, n822);
  and eco224 (patchNew_new_n400_, n953, patchNew_n1188);
  and eco225 (patchNew_new_n274_, n174, patchNew__not_GATE_23);
  and eco226 (patchNew_new_n265_, patchNew_new_n226_, patchNew__not_GATE_17);
  nor eco227 (patchNew_new_n377_, patchNew_new_n373_, patchNew_new_n376_);
  nor eco228 (patchNew_new_n431_, patchNew_new_n429_, patchNew_new_n430_);
  and eco229 (patchNew_new_n357_, patchNew_new_n353_, patchNew__not_GATE_53);
  nor eco230 (patchNew_new_n457_, n1168, patchNew_new_n455_);
  and eco231 (patchNew_new_n351_, patchNew_n1576, patchNew_n1584);
  and eco232 (patchNew_new_n370_, n793, patchNew__not_GATE_58);
  nor eco233 (patchNew_new_n446_, patchNew_new_n444_, patchNew_new_n445_);
  and eco234 (patchNew_new_n231_, patchNew__not_GATE_1, patchNew_new_n230_);
  and eco235 (patchNew_new_n297_, patchNew__not_GATE_33, patchNew_new_n296_);
  not eco236 (patchNew__not_GATE_71, n941);
  nor eco237 (patchNew_new_n257_, n587, patchNew_new_n255_);
  not eco238 (patchNew__not_GATE_2, patchNew_new_n231_);
  not eco239 (patchNew__not_GATE_85, n951);
  not eco240 (patchNew__not_GATE_3, n530);
  and eco241 (patchNew_new_n267_, patchNew__not_GATE_19, patchNew_new_n266_);
  not eco242 (patchNew__not_GATE_59, n793);
  and eco243 (patchNew_new_n308_, n1407, patchNew__xor_GATE_1);
  not eco244 (patchNew__not_GATE_55, patchNew_new_n358_);
  and eco245 (patchNew_new_n448_, n1147, patchNew_n1458);
  and eco246 (patchNew_new_n354_, n761, n727);
  nor eco247 (patchNew_new_n485_, patchNew_new_n447_, patchNew_new_n484_);
  nor eco248 (patchNew_new_n349_, patchNew_n1972, patchNew_new_n348_);
  and eco249 (patchNew_new_n295_, n17, n25);
  not eco250 (patchNew__not_GATE_4, patchNew_new_n235_);
  nor eco251 (patchNew_new_n480_, patchNew_new_n456_, patchNew_new_n479_);
  and eco252 (patchNew_new_n260_, patchNew__not_GATE_14, patchNew_new_n259_);
  not eco253 (patchNew__not_GATE_11, patchNew_new_n254_);
  and eco254 (patchNew_new_n302_, patchNew_new_n298_, patchNew_new_n301_);
  and eco255 (patchNew_new_n471_, patchNew_new_n454_, patchNew__xnor_GATE_9);
  nor eco256 (patchNew_new_n476_, n1204, patchNew_new_n455_);
  and eco257 (patchNew_new_n449_, n1115, n1131);
  and eco258 (patchNew_new_n411_, n935, patchNew__not_GATE_73);
  nor eco259 (patchNew_new_n253_, patchNew_new_n248_, patchNew_new_n251_);
  nor eco260 (patchNew_new_n363_, n713, patchNew_new_n362_);
  nor eco261 (patchNew_new_n375_, patchNew_new_n367_, patchNew_new_n374_);
  and eco262 (patchNew_new_n278_, n511, n624);
  not eco263 (patchNew__not_GATE_46, patchNew_new_n332_);
  and eco264 (patchNew_new_n290_, n1336, n1375);
  and eco265 (patchNew_new_n395_, n906, n890);
  not eco266 (patchNew__not_GATE_10, patchNew_n499);
  not eco267 (patchNew__not_GATE_56, patchNew_new_n360_);
  and eco268 (patchNew_new_n487_, patchNew__not_GATE_97, patchNew_new_n486_);
  nor eco269 (patchNew_new_n483_, patchNew_new_n423_, patchNew_new_n482_);
  nor eco270 (patchNew_new_n317_, patchNew_new_n315_, patchNew_new_n316_);
  not eco271 (patchNew__not_GATE_25, n1574);
  and eco272 (patchNew_new_n426_, patchNew_new_n422_, patchNew_new_n425_);
  and eco273 (patchNew_new_n232_, n638, patchNew__not_GATE_2);
  and eco274 (patchNew_new_n355_, patchNew__not_GATE_52, patchNew_n1384);
  and eco275 (patchNew_new_n493_, patchNew__not_GATE_100, patchNew_new_n492_);
  and eco276 (patchNew_new_n429_, patchNew__not_GATE_79, patchNew_new_n409_);
  and eco277 (patchNew_new_n437_, patchNew_new_n431_, patchNew__not_GATE_81);
  nor eco278 (patchNew_new_n532_, patchNew_new_n530_, patchNew_new_n531_);
  not eco279 (patchNew__not_GATE_114, n1546);
  not eco280 (patchNew__not_GATE_76, n1011);
  not eco281 (patchNew__not_GATE_43, patchNew_new_n302_);
  not eco282 (patchNew__not_GATE_94, patchNew_new_n475_);
  not eco283 (patchNew__not_GATE_62, n774);
  not eco284 (patchNew__not_GATE_84, n1012);
  and eco285 (patchNew_new_n416_, patchNew_new_n398_, patchNew__xnor_GATE_12);
  nor eco286 (patchNew_new_n417_, patchNew_new_n398_, patchNew__xnor_GATE_12);
  and eco287 (patchNew_new_n233_, patchNew__not_GATE_3, patchNew_n487);
  and eco288 (patchNew_new_n498_, patchNew_new_n349_, patchNew__xnor_GATE_7);
  nor eco289 (patchNew_new_n425_, patchNew_new_n410_, patchNew_new_n424_);
  and eco290 (patchNew_new_n303_, n586, patchNew__not_GATE_34);
  nor eco291 (patchNew_new_n465_, patchNew_new_n460_, patchNew_new_n463_);
  and eco292 (patchNew_new_n509_, patchNew_new_n428_, patchNew__not_GATE_105);
  and eco293 (patchNew_new_n407_, patchNew__not_GATE_71, patchNew_new_n406_);
  and eco294 (patchNew_new_n247_, patchNew__not_GATE_8, patchNew_new_n238_);
  nor eco295 (patchNew_new_n282_, n376, patchNew_new_n281_);
  nor eco296 (patchNew_new_n467_, n1193, patchNew_new_n466_);
  not eco297 (patchNew__not_GATE_27, patchNew_new_n282_);
  and eco298 (patchNew_new_n316_, n1962, patchNew_n844);
  and eco299 (patchNew_new_n423_, patchNew__not_GATE_78, patchNew_new_n422_);
  and eco300 (patchNew_new_n368_, patchNew__not_GATE_57, patchNew_new_n356_);
  and eco301 (patchNew_new_n475_, n1154, patchNew_new_n454_);
  nor eco302 (patchNew_new_n353_, patchNew_new_n351_, patchNew_new_n352_);
  not eco303 (patchNew__not_GATE_58, patchNew_new_n369_);
  nor eco304 (patchNew_new_n549_, patchNew_new_n547_, patchNew_new_n548_);
  nor eco305 (patchNew_new_n550_, patchNew_new_n489_, patchNew_new_n547_);
  and eco306 (patchNew_new_n234_, patchNew_n486, n478);
  nor eco307 (patchNew_new_n404_, patchNew_new_n398_, patchNew_new_n402_);
  not eco308 (patchNew__not_GATE_18, patchNew_n1020);
  nor eco309 (patchNew_new_n422_, patchNew_new_n419_, patchNew_new_n421_);
  not eco310 (patchNew__not_GATE_23, patchNew_new_n273_);
  nor eco311 (patchNew_new_n428_, patchNew_new_n426_, patchNew_new_n427_);
  nor eco312 (patchNew_new_n268_, patchNew_new_n232_, patchNew_new_n267_);
  and eco313 (patchNew_new_n405_, patchNew__not_GATE_70, patchNew_new_n404_);
  and eco314 (patchNew_new_n300_, n444, patchNew_new_n279_);
  nor eco315 (patchNew_new_n427_, patchNew_new_n422_, patchNew_new_n425_);
  nor eco316 (patchNew_new_n367_, patchNew_new_n361_, patchNew_new_n366_);
  not eco317 (patchNew__not_GATE_78, patchNew_new_n412_);
  and eco318 (patchNew_new_n430_, n928, patchNew_new_n406_);
  nor eco319 (patchNew_new_n238_, patchNew_new_n233_, patchNew_new_n237_);
  not eco320 (patchNew__not_GATE_63, patchNew_new_n384_);
  and eco321 (patchNew_new_n330_, patchNew__not_GATE_45, patchNew_new_n329_);
  nor eco322 (patchNew_new_n288_, n376, patchNew_new_n281_);
  nor eco323 (patchNew_new_n435_, patchNew_new_n388_, patchNew_new_n433_);
  and eco324 (patchNew_new_n391_, patchNew__not_GATE_66, patchNew_new_n390_);
  and eco325 (patchNew_new_n269_, patchNew__not_GATE_20, patchNew_new_n268_);
  not eco326 (patchNew__not_GATE_69, n854);
  not eco327 (patchNew__not_GATE_98, patchNew_new_n488_);
  nor eco328 (patchNew_new_n540_, patchNew_new_n274_, patchNew_new_n539_);
  and eco329 (patchNew_new_n541_, n138, patchNew__not_GATE_117);
  nor eco330 (patchNew_new_n589_, patchNew_new_n587_, patchNew_new_n588_);
  nor eco331 (patchNew_new_n590_, patchNew_new_n585_, patchNew_new_n589_);
  nor eco332 (patchNew_new_n591_, patchNew_new_n590_, patchNew__xor_GATE_1);
  and eco333 (patchNew_new_n481_, n1095, patchNew__not_GATE_96);
  and eco334 (patchNew_new_n266_, patchNew__not_GATE_18, n625);
  nor eco335 (patchNew_new_n454_, patchNew_new_n451_, patchNew_new_n453_);
  nor eco336 (patchNew_new_n358_, patchNew_new_n351_, patchNew_new_n357_);
  nor eco337 (patchNew_new_n286_, patchNew_new_n284_, patchNew_new_n285_);
  and eco338 (patchNew_new_n240_, n541, patchNew__not_GATE_5);
  nor eco339 (patchNew_new_n372_, patchNew_new_n370_, patchNew_new_n371_);
  not eco340 (patchNew__not_GATE_1, patchNew_new_n228_);
  not eco341 (patchNew__not_GATE_91, patchNew_n1469);
  not eco342 (patchNew__not_GATE_87, patchNew_new_n452_);
  not eco343 (patchNew__not_GATE_53, patchNew_new_n356_);
  nor eco344 (patchNew_new_n319_, patchNew_new_n308_, patchNew_new_n318_);
  nor eco345 (patchNew_new_n445_, patchNew_new_n418_, patchNew_new_n443_);
  and eco346 (patchNew_new_n474_, patchNew_new_n467_, patchNew_new_n473_);
  not eco347 (patchNew__not_GATE_34, patchNew_new_n255_);
  nor eco348 (patchNew_new_n436_, patchNew_new_n434_, patchNew_new_n435_);
  and eco349 (patchNew_new_n456_, n1168, patchNew_new_n455_);
  and eco350 (patchNew_new_n226_, n630, n634);
  not eco351 (patchNew__not_GATE_45, patchNew_new_n326_);
  nor eco352 (patchNew_new_n473_, patchNew_new_n471_, patchNew_new_n472_);
  nor eco353 (patchNew_new_n374_, patchNew_new_n370_, patchNew_new_n373_);
  not eco354 (patchNew__not_GATE_28, patchNew_new_n283_);
  and eco355 (patchNew_new_n547_, patchNew__not_GATE_120, patchNew_new_n546_);
  and eco356 (patchNew_new_n548_, patchNew_new_n545_, patchNew__not_GATE_121);
  and eco357 (patchNew_new_n244_, n613, patchNew_new_n243_);
  not eco358 (patchNew__not_GATE_7, n589);
  not eco359 (patchNew__not_GATE_42, patchNew_new_n321_);
  nor eco360 (patchNew_new_n482_, patchNew_new_n480_, patchNew_new_n481_);
  and eco361 (patchNew_new_n564_, patchNew_new_n510_, patchNew__not_GATE_128);
  not eco362 (patchNew__not_GATE_128, patchNew_new_n563_);
  not eco363 (patchNew__not_GATE_24, n174);
  nor eco364 (patchNew_new_n348_, patchNew_n1949, patchNew_new_n346_);
  nor eco365 (patchNew_new_n451_, n1106, patchNew_new_n450_);
  not eco366 (patchNew__not_GATE_57, patchNew_new_n353_);
  nor eco367 (patchNew_new_n466_, patchNew_new_n464_, patchNew_new_n465_);
  and eco368 (patchNew_new_n522_, patchNew__not_GATE_110, patchNew__xnor_GATE_8);
  not eco369 (patchNew__not_GATE_110, n1897);
  and eco370 (patchNew_new_n366_, patchNew_new_n358_, patchNew__not_GATE_56);
  not eco371 (patchNew__not_GATE_64, patchNew_new_n386_);
  nor eco372 (patchNew_new_n424_, n887, patchNew_new_n409_);
  xnor eco373 (patchNew__xnor_GATE_8, patchNew_new_n480_, patchNew_new_n518_);
  xnor eco374 (patchNew__xnor_GATE_9, n1154, n1204);
  xnor eco375 (patchNew__xnor_GATE_10, patchNew_new_n319_, patchNew_new_n323_);
  xnor eco376 (patchNew__xnor_GATE_11, patchNew_new_n504_, patchNew_new_n510_);
  xnor eco377 (patchNew__xnor_GATE_12, n953, n952);
  xnor eco378 (patchNew__xnor_GATE_13, patchNew_new_n556_, patchNew_new_n557_);
  nor eco379 (patchNew_new_n499_, patchNew_new_n349_, patchNew__xnor_GATE_7);
  and eco380 (patchNew_new_n501_, patchNew_new_n325_, patchNew_new_n329_);
  not eco381 (patchNew__not_GATE_88, patchNew_new_n454_);
  nor eco382 (patchNew_new_n576_, patchNew_new_n574_, patchNew_new_n575_);
  not eco383 (patchNew__not_GATE_131, patchNew_new_n570_);
  and eco384 (patchNew_new_n236_, n514, patchNew__not_GATE_4);
  and eco385 (patchNew_new_n599_, n1666, patchNew_new_n323_);
  nor eco386 (patchNew_new_n600_, patchNew_new_n529_, patchNew_new_n599_);
  nor eco387 (patchNew_new_n601_, patchNew_new_n597_, patchNew_new_n600_);
  and eco388 (patchNew_new_n602_, patchNew__not_GATE_141, patchNew_new_n601_);
  and eco389 (patchNew_new_n536_, patchNew_new_n532_, patchNew__xnor_GATE_10);
  nor eco390 (patchNew_new_n325_, patchNew_new_n320_, patchNew_new_n324_);
  not eco391 (patchNew__not_GATE_103, patchNew_new_n446_);
  nor eco392 (patchNew_new_n510_, patchNew_new_n508_, patchNew_new_n509_);
  and eco393 (patchNew_new_n572_, patchNew__not_GATE_132, patchNew_new_n570_);
  not eco394 (patchNew__not_GATE_132, n1710);
  and eco395 (patchNew_new_n565_, patchNew__not_GATE_129, patchNew__xor_GATE_1);
  not eco396 (patchNew__not_GATE_129, n1754);
  nor eco397 (patchNew_new_n619_, n1614, patchNew_new_n618_);
  and eco398 (patchNew_new_n620_, patchNew__not_GATE_150, patchNew_new_n618_);
  not eco399 (patchNew__not_GATE_150, n674);
  nor eco400 (patchNew_new_n621_, patchNew_new_n619_, patchNew_new_n620_);
  and eco401 (patchNew_new_n622_, patchNew__not_GATE_151, patchNew_new_n621_);
  nor eco402 (patchNew_new_n323_, patchNew_new_n262_, patchNew_new_n322_);
  not eco403 (patchNew__not_GATE_19, patchNew_new_n265_);
  nor eco404 (patchNew_new_n259_, patchNew_new_n243_, patchNew_new_n258_);
  and eco405 (patchNew_new_n270_, n642, patchNew__not_GATE_21);
  and eco406 (patchNew_new_n310_, patchNew__not_GATE_37, patchNew_new_n254_);
  and eco407 (patchNew_new_n464_, patchNew_new_n460_, patchNew_new_n463_);
  nor eco408 (patchNew_new_n678_, patchNew_new_n593_, patchNew_new_n677_);
  and eco409 (patchNew_new_n680_, n1754, n1699);
  and eco410 (patchNew_new_n681_, patchNew_new_n590_, patchNew__not_GATE_167);
  not eco411 (patchNew__not_GATE_167, patchNew_new_n680_);
  nor eco412 (patchNew_new_n682_, patchNew_new_n583_, patchNew_new_n587_);
  nor eco413 (patchNew_new_n329_, patchNew_new_n327_, patchNew_new_n328_);
  nor eco414 (patchNew_new_n412_, patchNew_new_n410_, patchNew_new_n411_);
  and eco415 (patchNew_new_n410_, n887, patchNew_new_n409_);
  nor eco416 (patchNew_new_n420_, n1012, patchNew_new_n418_);
  and eco417 (patchNew_new_n333_, n1381, patchNew__not_GATE_46);
  not eco418 (patchNew__not_GATE_121, patchNew_new_n546_);
  not eco419 (patchNew__not_GATE_118, n138);
  and eco420 (patchNew_new_n440_, patchNew__not_GATE_83, patchNew_new_n436_);
  not eco421 (patchNew__not_GATE_14, patchNew_new_n257_);
  nor eco422 (patchNew_new_n409_, patchNew_new_n407_, patchNew_new_n408_);
  and eco423 (patchNew_new_n442_, patchNew__not_GATE_85, n1012);
  and eco424 (patchNew_new_n586_, n1193, patchNew_new_n466_);
  and eco425 (patchNew_new_n582_, n1754, n1708);
  nor eco426 (patchNew_new_n583_, patchNew_new_n581_, patchNew_new_n582_);
  and eco427 (patchNew_new_n544_, patchNew_new_n393_, patchNew__not_GATE_119);
  nor eco428 (patchNew_new_n545_, patchNew_new_n391_, patchNew_new_n544_);
  nor eco429 (patchNew_new_n460_, patchNew_new_n452_, patchNew_new_n459_);
  and eco430 (patchNew_new_n227_, n378, n439);
  not eco431 (patchNew__not_GATE_54, patchNew_n1642);
  and eco432 (patchNew_new_n462_, patchNew__not_GATE_91, n1070);
  not eco433 (patchNew__not_GATE_26, patchNew_new_n280_);
  not eco434 (patchNew__not_GATE_72, patchNew_new_n406_);
  not eco435 (patchNew__not_GATE_65, patchNew_new_n379_);
  and eco436 (patchNew_new_n479_, patchNew_new_n458_, patchNew__not_GATE_95);
  and eco437 (patchNew_new_n328_, n512, patchNew_new_n263_);
  not eco438 (patchNew__not_GATE_151, patchNew_new_n615_);
  nor eco439 (patchNew_new_n623_, patchNew_new_n621_, patchNew__xnor_GATE_7);
  and eco440 (patchNew_new_n624_, patchNew_new_n554_, patchNew_new_n623_);
  nor eco441 (patchNew_new_n625_, patchNew_new_n622_, patchNew_new_n624_);
  xnor eco442 (patchNew__xnor_GATE_0, patchNew_new_n517_, patchNew_new_n524_);
  xor eco443 (patchNew__xor_GATE_1, patchNew_new_n304_, patchNew_new_n259_);
  and eco444 (patchNew_new_n687_, patchNew__not_GATE_170, patchNew_new_n680_);
  not eco445 (patchNew__not_GATE_170, patchNew_new_n576_);
  and eco446 (patchNew_new_n688_, patchNew_new_n583_, patchNew__not_GATE_171);
  and eco447 (patchNew_new_n690_, n1666, n2007);
  not eco448 (patchNew__not_GATE_171, patchNew_new_n687_);
  and eco449 (patchNew_new_n542_, patchNew__not_GATE_118, patchNew_new_n540_);
  and eco450 (patchNew_new_n611_, patchNew_new_n610_, patchNew__xnor_GATE_13);
  and eco451 (patchNew_new_n612_, patchNew__not_GATE_147, patchNew_new_n487_);
  not eco452 (patchNew__not_GATE_147, patchNew_new_n393_);
  and eco453 (patchNew_new_n492_, patchNew_new_n365_, patchNew__not_GATE_99);
  nor eco454 (patchNew_new_n332_, patchNew_new_n302_, patchNew_new_n331_);
  not eco455 (patchNew__not_GATE_99, patchNew_new_n375_);
  nor eco456 (patchNew_new_n293_, n17, n25);
  and eco457 (patchNew_new_n239_, n540, patchNew_new_n238_);
  not eco458 (patchNew__not_GATE_95, patchNew_new_n478_);
  and eco459 (patchNew_new_n346_, patchNew_new_n342_, patchNew__xnor_GATE_3);
  nor eco460 (patchNew_new_n566_, patchNew_new_n467_, patchNew_new_n473_);
  nor eco461 (patchNew_new_n567_, patchNew_new_n474_, patchNew_new_n566_);
  nor eco462 (patchNew_new_n568_, patchNew_new_n565_, patchNew_new_n567_);
  not eco463 (patchNew__not_GATE_144, patchNew_new_n329_);
  and eco464 (patchNew_new_n607_, patchNew__not_GATE_145, patchNew_new_n606_);
  not eco465 (patchNew__not_GATE_145, patchNew_new_n605_);
  and eco466 (patchNew_new_n408_, n941, patchNew__not_GATE_72);
  nor eco467 (patchNew_new_n478_, patchNew_new_n474_, patchNew_new_n477_);
  xnor eco468 (patchNew__xnor_GATE_2, patchNew_new_n550_, patchNew_new_n365_);
  xnor eco469 (patchNew__xnor_GATE_3, n211, patchNew_new_n270_);
  not eco470 (patchNew__not_GATE_68, patchNew_new_n401_);
  nor eco471 (patchNew_new_n598_, patchNew_new_n529_, patchNew_new_n595_);
  nor eco472 (patchNew_new_n587_, patchNew_new_n467_, patchNew_new_n586_);
  nor eco473 (patchNew_new_n588_, patchNew_n844, patchNew_new_n577_);
  and eco474 (patchNew_new_n604_, patchNew__not_GATE_143, patchNew__xnor_GATE_8);
  not eco475 (patchNew__not_GATE_143, patchNew_new_n603_);
  nor eco476 (patchNew_new_n605_, patchNew_new_n602_, patchNew__xnor_GATE_8);
  and eco477 (patchNew_new_n606_, n1666, patchNew__not_GATE_144);
  nor eco478 (patchNew_new_n502_, n1897, patchNew_new_n331_);
  nor eco479 (patchNew_new_n503_, patchNew_new_n501_, patchNew_new_n502_);
  nor eco480 (patchNew_new_n506_, patchNew_new_n480_, patchNew_new_n505_);
  nor eco481 (patchNew_new_n507_, patchNew_new_n447_, patchNew_new_n506_);
  and eco482 (patchNew_new_n554_, patchNew_new_n549_, patchNew__xnor_GATE_2);
  and eco483 (patchNew_new_n555_, patchNew_new_n544_, patchNew_new_n554_);
  and eco484 (patchNew_new_n283_, n634, patchNew__not_GATE_27);
  and eco485 (patchNew_new_n514_, patchNew_new_n503_, patchNew__xnor_GATE_11);
  nor eco486 (patchNew_new_n515_, patchNew_new_n503_, patchNew__xnor_GATE_11);
  nor eco487 (patchNew_new_n613_, patchNew_new_n611_, patchNew_new_n612_);
  nor eco488 (patchNew_new_n614_, patchNew_new_n555_, patchNew_new_n613_);
  and eco489 (patchNew_new_n615_, patchNew__not_GATE_148, patchNew_new_n614_);
  not eco490 (patchNew__not_GATE_148, patchNew__xnor_GATE_7);
  not eco491 (patchNew__not_GATE_120, patchNew_new_n545_);
  and eco492 (patchNew_new_n419_, patchNew__not_GATE_76, patchNew_new_n418_);
  not eco493 (patchNew__not_GATE_90, n1070);
  nor eco494 (patchNew_new_n543_, patchNew_new_n541_, patchNew_new_n542_);
  not eco495 (patchNew__not_GATE_117, patchNew_new_n540_);
  nor eco496 (patchNew_new_n556_, patchNew_new_n437_, patchNew_new_n440_);
  nor eco497 (patchNew_new_n557_, patchNew_new_n423_, patchNew_new_n509_);
  nor eco498 (patchNew_new_n401_, patchNew_new_n399_, patchNew_new_n400_);
  not eco499 (patchNew__not_GATE_89, patchNew_new_n450_);
  nor eco500 (patchNew_new_n546_, patchNew_new_n375_, patchNew_new_n489_);
  not eco501 (patchNew__not_GATE_119, patchNew_new_n487_);
  nor eco502 (patchNew_new_n418_, patchNew_new_n416_, patchNew_new_n417_);
  nor eco503 (patchNew_new_n584_, patchNew_n844, patchNew_new_n583_);
  and eco504 (patchNew_new_n585_, n1666, patchNew__not_GATE_138);
  not eco505 (patchNew__not_GATE_138, patchNew_new_n584_);
  nor eco506 (patchNew_new_n517_, patchNew_new_n331_, patchNew_new_n501_);
  nor eco507 (patchNew_new_n518_, patchNew_new_n447_, patchNew_new_n481_);
  and eco508 (patchNew_new_n488_, patchNew_new_n393_, patchNew_new_n487_);
  and eco509 (patchNew_new_n388_, patchNew__not_GATE_64, patchNew_new_n387_);
  and eco510 (patchNew_new_n235_, n477, n535);
  and eco511 (patchNew_new_n285_, n331, patchNew_new_n283_);
  not eco512 (patchNew__not_GATE_16, patchNew_new_n263_);
  nor eco513 (patchNew_new_n581_, patchNew_new_n577_, patchNew_new_n580_);
  and eco514 (patchNew_new_n580_, n1454, patchNew__not_GATE_137);
  not eco515 (patchNew__not_GATE_137, patchNew_new_n579_);
  and eco516 (patchNew_new_n461_, patchNew_n1469, patchNew__not_GATE_90);
  and eco517 (patchNew_new_n229_, n334, n374);
  not eco518 (patchNew__not_GATE_5, patchNew_new_n238_);
  and eco519 (patchNew_new_n322_, patchNew__not_GATE_41, patchNew_new_n261_);
  and eco520 (patchNew_new_n638_, patchNew__not_GATE_155, patchNew_n1720);
  not eco521 (patchNew__not_GATE_149, patchNew_new_n494_);
  and eco522 (patchNew_new_n617_, patchNew_n1705, patchNew_n1706);
  nor eco523 (patchNew_new_n618_, patchNew_new_n616_, patchNew_new_n617_);
  nor eco524 (patchNew_new_n369_, patchNew_new_n357_, patchNew_new_n368_);
  and eco525 (patchNew_new_n575_, n1754, patchNew__not_GATE_135);
  nor eco526 (patchNew_new_n579_, n1708, patchNew_new_n578_);
  not eco527 (patchNew__not_GATE_135, patchNew_new_n571_);
  nor eco528 (patchNew_new_n651_, patchNew_new_n549_, patchNew_n1911);
  and eco529 (patchNew_new_n653_, patchNew_n1063, patchNew_new_n549_);
  nor eco530 (patchNew_new_n654_, patchNew_n1063, patchNew_new_n549_);
  and eco531 (patchNew_new_n656_, patchNew__not_GATE_159, patchNew_n1907);
  not eco532 (patchNew__not_GATE_159, patchNew_new_n611_);
  and eco533 (patchNew_new_n670_, n1754, patchNew_new_n567_);
  not eco534 (patchNew__not_GATE_160, patchNew_new_n286_);
  and eco535 (patchNew_new_n577_, n1708, patchNew_new_n576_);
  and eco536 (patchNew_new_n578_, n1666, patchNew__not_GATE_136);
  not eco537 (patchNew__not_GATE_136, patchNew_new_n574_);
  not eco538 (patchNew__not_GATE_155, patchNew_new_n623_);
  not eco539 (patchNew__not_GATE_156, patchNew_new_n635_);
  nor eco540 (patchNew_new_n640_, n137, n136);
  and eco541 (patchNew_new_n641_, n138, patchNew__not_GATE_157);
  not eco542 (patchNew__not_GATE_157, patchNew_new_n540_);
  not eco543 (patchNew__not_GATE_113, patchNew_new_n458_);
  nor eco544 (patchNew_new_n529_, patchNew_new_n479_, patchNew_new_n528_);
  and eco545 (patchNew_new_n563_, n1666, patchNew__not_GATE_127);
  not eco546 (patchNew__not_GATE_127, patchNew_new_n301_);
  not eco547 (patchNew__not_GATE_153, patchNew_new_n337_);
  nor eco548 (patchNew_new_n635_, patchNew_new_n614_, patchNew__xnor_GATE_7);
  nor eco549 (patchNew_new_n636_, n1614, patchNew_new_n618_);
  nor eco550 (patchNew_new_n658_, patchNew_new_n610_, patchNew__xnor_GATE_13);
  not eco551 (patchNew__not_GATE_154, patchNew_new_n636_);
  not eco552 (patchNew__not_GATE_73, patchNew_new_n409_);
  nor eco553 (patchNew_new_n390_, patchNew_new_n378_, patchNew_new_n389_);
  and eco554 (patchNew_new_n477_, patchNew__not_GATE_94, patchNew_new_n476_);
  nor eco555 (patchNew_new_n523_, n1381, patchNew__xnor_GATE_8);
  and eco556 (patchNew_new_n389_, patchNew__not_GATE_65, patchNew_new_n388_);
  xnor eco557 (patchNew__xnor_GATE_4, patchNew_new_n317_, patchNew_new_n567_);
  xnor eco558 (patchNew__xnor_GATE_5, n1424, patchNew_new_n587_);
  xnor eco559 (patchNew__xnor_GATE_6, patchNew_new_n621_, patchNew_new_n543_);
  xnor eco560 (patchNew__xnor_GATE_7, n1778, patchNew_new_n494_);
  and eco561 (patchNew_new_n561_, patchNew__not_GATE_126, patchNew_new_n301_);
  and eco562 (patchNew_new_n528_, patchNew__not_GATE_113, patchNew_new_n478_);
  not eco563 (patchNew__not_GATE_100, patchNew_new_n491_);
  not eco564 (patchNew__not_GATE_83, patchNew_new_n431_);
  not eco565 (patchNew__not_GATE_133, n1461);
  and eco566 (patchNew_new_n574_, patchNew__not_GATE_134, patchNew_n1791);
  not eco567 (patchNew__not_GATE_134, patchNew_new_n571_);
  and eco568 (patchNew_new_n327_, n1386, patchNew__not_GATE_44);
  and eco569 (patchNew_new_n455_, n1206, patchNew__not_GATE_88);
  nor eco570 (patchNew_new_n524_, patchNew_new_n522_, patchNew_new_n523_);
  nor eco571 (patchNew_new_n486_, patchNew_new_n439_, patchNew_new_n440_);
  and eco572 (patchNew_new_n571_, n1710, patchNew__not_GATE_131);
  not eco573 (patchNew__not_GATE_126, n1754);
  nor eco574 (patchNew_new_n490_, patchNew_new_n391_, patchNew_new_n489_);
  and eco575 (patchNew_new_n491_, patchNew__not_GATE_98, patchNew_new_n490_);
  not eco576 (patchNew__not_GATE_141, patchNew_new_n598_);
  and eco577 (patchNew_new_n603_, n1666, patchNew__not_GATE_142);
  not eco578 (patchNew__not_GATE_142, patchNew_new_n602_);
  and eco579 (patchNew_new_n569_, n1627, n1718);
  and eco580 (patchNew_new_n570_, n1717, patchNew__not_GATE_130);
  not eco581 (patchNew__not_GATE_130, patchNew_new_n569_);
  nor eco582 (patchNew_new_n331_, patchNew_new_n325_, patchNew_new_n329_);
  not eco583 (patchNew__not_GATE_66, patchNew_new_n377_);
  and eco584 (patchNew_new_n597_, patchNew__not_GATE_140, patchNew_new_n596_);
  nor eco585 (patchNew_new_n610_, patchNew_new_n562_, patchNew_new_n609_);
  not eco586 (patchNew__not_GATE_140, patchNew_new_n595_);
  nor eco587 (patchNew_new_n594_, patchNew_new_n567_, patchNew_new_n590_);
  nor eco588 (patchNew_new_n595_, patchNew_new_n593_, patchNew_new_n594_);
  nor eco589 (patchNew_new_n596_, n1754, patchNew_new_n323_);
  and eco590 (patchNew_new_n392_, patchNew_new_n377_, patchNew__not_GATE_67);
  nor eco591 (patchNew_new_n562_, patchNew_new_n510_, patchNew_new_n561_);
  and eco592 (patchNew_new_n508_, patchNew__not_GATE_104, patchNew_new_n507_);
  not eco593 (patchNew__not_GATE_104, patchNew_new_n428_);
  and eco594 (patchNew_new_n643_, patchNew_new_n614_, patchNew__xnor_GATE_7);
  and eco595 (patchNew_new_n645_, n1597, patchNew_new_n540_);
  and eco596 (patchNew_new_n646_, patchNew_n1972, patchNew__not_GATE_158);
  not eco597 (patchNew__not_GATE_158, patchNew_new_n645_);
  and eco598 (patchNew_new_n648_, patchNew_new_n549_, patchNew_n1911);
  nor eco599 (patchNew_new_n649_, patchNew_new_n648_, patchNew__xnor_GATE_2);
  and eco600 (patchNew_new_n326_, patchNew__not_GATE_43, patchNew_new_n325_);
  nor eco601 (patchNew_new_n626_, patchNew_new_n543_, patchNew_new_n625_);
  not eco602 (patchNew__not_GATE_152, patchNew_n1907);
  nor eco603 (patchNew_new_n629_, patchNew_new_n621_, patchNew_n1911);
  nor eco604 (patchNew_new_n631_, patchNew_new_n342_, patchNew__xnor_GATE_3);
  and eco605 (patchNew_new_n633_, patchNew_new_n286_, patchNew__not_GATE_153);
  and eco606 (patchNew_new_n592_, n1666, patchNew__not_GATE_139);
  not eco607 (patchNew__not_GATE_139, patchNew_new_n591_);
  nor eco608 (patchNew_new_n593_, patchNew_new_n568_, patchNew_new_n592_);
  and eco609 (patchNew_new_n530_, patchNew__not_GATE_114, patchNew_new_n529_);
  nor eco610 (patchNew_new_n531_, n1555, patchNew_new_n529_);
  not eco611 (patchNew__not_GATE_0, patchNew_new_n229_);
  nor eco612 (patchNew_new_n494_, patchNew_new_n363_, patchNew_new_n493_);
  nor eco613 (patchNew_new_n365_, patchNew_new_n363_, patchNew_new_n364_);
  not eco614 (patchNew__not_GATE_67, patchNew_new_n390_);
  and eco615 (patchNew_new_n258_, n589, patchNew__not_GATE_13);
  nor eco616 (patchNew_new_n537_, patchNew_new_n532_, patchNew__xnor_GATE_10);
  and eco617 (patchNew_new_n539_, patchNew_n1047, patchNew_n1050);
  and eco618 (patchNew_new_n324_, patchNew__not_GATE_42, patchNew_new_n323_);
  not eco619 (patchNew__not_GATE_44, patchNew_new_n263_);
  and eco620 (patchNew_new_n403_, patchNew__not_GATE_69, patchNew_new_n401_);
  and eco621 (patchNew_new_n660_, n1754, patchNew__xnor_GATE_8);
  not eco622 (patchNew__not_GATE_161, patchNew_new_n660_);
  and eco623 (patchNew_new_n662_, patchNew__not_GATE_162, patchNew_new_n608_);
  not eco624 (patchNew__not_GATE_162, patchNew_new_n510_);
  and eco625 (patchNew_new_n664_, patchNew_n1989, patchNew__xnor_GATE_13);
  nor eco626 (patchNew_new_n665_, patchNew_n1989, patchNew__xnor_GATE_13);
  and eco627 (patchNew_new_n667_, n1754, patchNew_new_n529_);
  not eco628 (patchNew__not_GATE_163, patchNew_new_n329_);
  nor eco629 (patchNew_new_n608_, patchNew_new_n604_, patchNew_new_n607_);
  and eco630 (patchNew_new_n609_, patchNew__not_GATE_146, patchNew_new_n608_);
  and eco631 (patchNew_new_n616_, n711, patchNew__not_GATE_149);
  not eco632 (patchNew__not_GATE_146, patchNew_new_n564_);
  and eco633 (patchNew_new_n505_, n1095, patchNew__not_GATE_103);
  and eco634 (patchNew_new_n489_, patchNew_new_n367_, patchNew_new_n374_);
  not eco635 (patchNew__not_GATE_164, patchNew_new_n670_);
  and eco636 (patchNew_new_n677_, n1754, patchNew_new_n587_);
  not eco637 (patchNew_n499, patchNew_n437);
  xor eco638 (patchNew_n1390, patchNew_n1367, patchNew_n1389);
  xnor eco639 (patchNew_n1224, patchNew_n1210, patchNew_n1223);
  nand eco640 (patchNew_n1008, patchNew_n996, patchNew_n1007);
  xor eco641 (patchNew_n989, patchNew_n986, n168);
  xor eco642 (patchNew_n1188, n846, n834);
  xnor eco643 (patchNew_n1576, patchNew_n1572, patchNew_n1575);
  xor eco644 (patchNew_n1584, patchNew_n1582, n692);
  xor eco645 (patchNew_n1458, patchNew_n1455, patchNew_n1457);
  xor eco646 (patchNew_n1384, patchNew_n1373, patchNew_n1383);
  xnor eco647 (patchNew_n487, patchNew_n484, patchNew_n486);
  nand eco648 (patchNew_n486, patchNew_n485, patchNew_n429);
  nor eco649 (patchNew_n1020, n330, n264);
  not eco650 (patchNew_n1469, patchNew_n1433);
  xnor eco651 (patchNew_n1642, patchNew_n1630, patchNew_n1641);
  nand eco652 (patchNew_n1705, patchNew_n1703, patchNew_n1704);
  xor eco653 (patchNew_n1706, n667, patchNew_n1100);
  xor eco654 (patchNew_n1047, patchNew_n951, patchNew_n952);
  nand eco655 (patchNew_n1050, patchNew_n1048, patchNew_n1049);
  xnor eco656 (patchNew_n437, patchNew_n435, patchNew_n436);
  nand eco657 (patchNew_n1367, patchNew_n1364, patchNew_n1366);
  or eco658 (patchNew_n1389, patchNew_n1385, patchNew_n1388);
  xor eco659 (patchNew_n1210, n867, n864);
  nor eco660 (patchNew_n1223, patchNew_n1221, patchNew_n1222);
  or eco661 (patchNew_n996, patchNew_n992, n207);
  nand eco662 (patchNew_n1007, patchNew_n1002, patchNew_n1006);
  xnor eco663 (patchNew_n986, n164, n165);
  xor eco664 (patchNew_n1572, n685, patchNew_n1376);
  nand eco665 (patchNew_n1575, patchNew_n1377, patchNew_n1574);
  nand eco666 (patchNew_n1582, patchNew_n1580, patchNew_n1581);
  xor eco667 (patchNew_n1455, n1056, n1115);
  nand eco668 (patchNew_n1457, patchNew_n1456, patchNew_n1422);
  xor eco669 (patchNew_n1373, n679, n761);
  nand eco670 (patchNew_n1383, patchNew_n1377, patchNew_n1382);
  xor eco671 (patchNew_n484, n476, n515);
  not eco672 (patchNew_n485, patchNew_n427);
  nand eco673 (patchNew_n429, n533, n479);
  xnor eco674 (patchNew_n1433, patchNew_n1430, patchNew_n1432);
  xor eco675 (patchNew_n1630, patchNew_n1627, n698);
  nand eco676 (patchNew_n1641, patchNew_n1638, patchNew_n1640);
  or eco677 (patchNew_n1703, n705, patchNew_n1702);
  or eco678 (patchNew_n1704, n701, n702);
  nor eco679 (patchNew_n1100, patchNew_n1098, patchNew_n1099);
  nor eco680 (patchNew_n951, patchNew_n948, patchNew_n950);
  not eco681 (patchNew_n952, n131);
  or eco682 (patchNew_n1048, patchNew_n986, n168);
  or eco683 (patchNew_n1049, n164, n165);
  xor eco684 (patchNew_n435, n473, n397);
  nand eco685 (patchNew_n436, patchNew_n375, patchNew_n370);
  or eco686 (patchNew_n1364, patchNew_n1354, n785);
  nand eco687 (patchNew_n1366, patchNew_n1365, n785);
  and eco688 (patchNew_n1385, n721, patchNew_n1384);
  and eco689 (patchNew_n1388, patchNew_n1386, patchNew_n1387);
  and eco690 (patchNew_n1221, n782, n762);
  and eco691 (patchNew_n1222, n781, n866);
  not eco692 (patchNew_n992, patchNew_n991);
  not eco693 (patchNew_n1002, patchNew_n1001);
  nand eco694 (patchNew_n1006, patchNew_n1003, patchNew_n1005);
  not eco695 (patchNew_n1376, n683);
  nand eco696 (patchNew_n1377, patchNew_n1374, patchNew_n1376);
  nand eco697 (patchNew_n1574, patchNew_n1573, patchNew_n1382);
  not eco698 (patchNew_n1580, n694);
  or eco699 (patchNew_n1581, n890, n673);
  not eco700 (patchNew_n1456, patchNew_n1425);
  nand eco701 (patchNew_n1422, n1059, n1126);
  nand eco702 (patchNew_n1382, n677, n676);
  nor eco703 (patchNew_n427, n533, n479);
  xor eco704 (patchNew_n1430, n1053, n1075);
  nand eco705 (patchNew_n1432, patchNew_n1431, patchNew_n1284);
  nor eco706 (patchNew_n1627, patchNew_n1626, n694);
  or eco707 (patchNew_n1638, patchNew_n1631, patchNew_n1637);
  nand eco708 (patchNew_n1640, patchNew_n1639, patchNew_n1575);
  not eco709 (patchNew_n1702, n712);
  and eco710 (patchNew_n1098, n666, patchNew_n1097);
  and eco711 (patchNew_n1099, patchNew_n1094, n669);
  and eco712 (patchNew_n948, patchNew_n945, patchNew_n947);
  and eco713 (patchNew_n950, n130, n133);
  nand eco714 (patchNew_n375, n487, n389);
  nand eco715 (patchNew_n370, n496, n407);
  not eco716 (patchNew_n1354, n790);
  not eco717 (patchNew_n1365, n790);
  not eco718 (patchNew_n1386, n721);
  not eco719 (patchNew_n1387, patchNew_n1384);
  not eco720 (patchNew_n991, n204);
  nor eco721 (patchNew_n1001, patchNew_n999, patchNew_n1000);
  or eco722 (patchNew_n1003, patchNew_n614, n195);
  or eco723 (patchNew_n1005, n200, n197);
  not eco724 (patchNew_n1374, n717);
  not eco725 (patchNew_n1573, n679);
  nor eco726 (patchNew_n1425, n1126, n1059);
  not eco727 (patchNew_n1431, patchNew_n1289);
  nand eco728 (patchNew_n1284, n1076, n1004);
  and eco729 (patchNew_n1626, patchNew_n1581, n692);
  not eco730 (patchNew_n1631, patchNew_n1376);
  not eco731 (patchNew_n1637, patchNew_n1636);
  not eco732 (patchNew_n1639, n685);
  not eco733 (patchNew_n1097, n669);
  nor eco734 (patchNew_n1094, patchNew_n1092, patchNew_n1093);
  nor eco735 (patchNew_n945, patchNew_n943, patchNew_n944);
  not eco736 (patchNew_n947, n133);
  and eco737 (patchNew_n999, n207, patchNew_n998);
  and eco738 (patchNew_n1000, patchNew_n994, n204);
  not eco739 (patchNew_n614, patchNew_n613);
  nor eco740 (patchNew_n1289, n891, n1066);
  nand eco741 (patchNew_n1636, patchNew_n1634, patchNew_n1635);
  and eco742 (patchNew_n1092, patchNew_n1091, n661);
  and eco743 (patchNew_n1093, n660, n663);
  and eco744 (patchNew_n943, patchNew_n942, n125);
  and eco745 (patchNew_n944, n124, n127);
  not eco746 (patchNew_n998, n204);
  xnor eco747 (patchNew_n994, patchNew_n993, patchNew_n971);
  nand eco748 (patchNew_n613, patchNew_n611, patchNew_n612);
  or eco749 (patchNew_n1634, patchNew_n1632, n682);
  or eco750 (patchNew_n1635, patchNew_n1575, n685);
  xor eco751 (patchNew_n1091, n660, n663);
  xor eco752 (patchNew_n942, n124, n127);
  xor eco753 (patchNew_n993, patchNew_n976, n161);
  nand eco754 (patchNew_n971, patchNew_n968, patchNew_n970);
  or eco755 (patchNew_n611, patchNew_n600, n200);
  or eco756 (patchNew_n612, patchNew_n609, n197);
  not eco757 (patchNew_n1632, n685);
  nor eco758 (patchNew_n976, patchNew_n975, n157);
  or eco759 (patchNew_n968, patchNew_n961, patchNew_n967);
  nand eco760 (patchNew_n970, patchNew_n969, patchNew_n608);
  not eco761 (patchNew_n600, n197);
  xnor eco762 (patchNew_n609, patchNew_n603, patchNew_n608);
  and eco763 (patchNew_n975, patchNew_n592, n155);
  not eco764 (patchNew_n961, patchNew_n602);
  not eco765 (patchNew_n967, patchNew_n966);
  not eco766 (patchNew_n969, n148);
  nand eco767 (patchNew_n608, patchNew_n606, patchNew_n607);
  xor eco768 (patchNew_n603, n148, patchNew_n602);
  or eco769 (patchNew_n592, n342, n137);
  not eco770 (patchNew_n602, n146);
  nand eco771 (patchNew_n966, patchNew_n964, patchNew_n965);
  or eco772 (patchNew_n606, n142, n144);
  not eco773 (patchNew_n607, patchNew_n201);
  or eco774 (patchNew_n964, patchNew_n962, n145);
  or eco775 (patchNew_n965, patchNew_n608, n148);
  nor eco776 (patchNew_n201, n146, n179);
  not eco777 (patchNew_n962, n148);
endmodule
