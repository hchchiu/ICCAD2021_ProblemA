module top_eco(\y[7]_in, \a[0], n_490, \op[0], \a[1], \a[2], \a[3], \a[4], \a[5], \b[0], \b[1], \b[2], \b[3], \b[4], \b[5], \op[1], n_505, n_506, wc1, n_474, wc3, n_482, n_489, wc7, n_565, n_571, wc17, wc20, n_508, wc21, wc22, n_665, wc52, wc26, n_492, wc27, n_713, n_668, wc42, n_472, wc47, n_471, n_710, n_582, n_725, n_680, n_695, wc61, overflow, \y[0], parity, \y[1], \y[2], \y[3], \y[4], \y[5], \y[6], \y[7]);
  input \y[7]_in, \a[0], n_490, \op[0], \a[1];
  input \a[2], \a[3], \a[4], \a[5], \b[0];
  input \b[1], \b[2], \b[3], \b[4], \b[5];
  input \op[1], n_505, n_506, wc1, n_474;
  input wc3, n_482, n_489, wc7, n_565;
  input n_571, wc17, wc20, n_508, wc21;
  input wc22, n_665, wc52, wc26, n_492;
  input wc27, n_713, n_668, wc42, n_472;
  input wc47, n_471, n_710, n_582, n_725;
  input n_680, n_695, wc61;
  output overflow, \y[0], parity, \y[1], \y[2];
  output \y[3], \y[4], \y[5], \y[6], \y[7];
  wire nn_539, nn_264, nn_475, nn_496, nn_535;
  wire nn_803, nn_540, nn_541, nn_802, nwc10;
  wire nn_195, nn_451, nwc28, nn_551, nn_804;
  wire nwc12, nn_450, nn_502, nn_805, nwc13;
  wire nn_806, nn_193, nn_190, nn_807, nwc16;
  wire nn_729, nn_728, nn_811, nn_140, nn_544;
  wire nwc17, nn_191, nn_503, nn_812, nn_726;
  wire nn_727, nn_69, nn_505, nwc19, nn_783;
  wire nn_782, nwc21, nn_545, nn_696, nwc23;
  wire nn_780, nn_701, nn_702, nn_550, nn_455;
  wire nn_705, nn_819, nn_820, nn_694, nn_695;
  wire nn_413, nn_185, nn_453, nn_670, nwc30;
  wire nwc31, nn_672, nwc32, nn_522, nn_671;
  wire nn_687, nn_683, nn_677, nn_678, nn_47;
  wire nwc34, nn_759, nn_758, nwc37, nn_369;
  wire nwc38, nn_410, nn_756, nn_552, nn_657;
  wire nn_662, nn_597, nwc41, nwc42, nn_553;
  wire nn_56, nn_611, nn_620, nn_602, nn_603;
  wire nn_595, nn_596, nn_521, nn_615, nn_41;
  wire nn_612, nwc48, nn_360, nwc49, nn_543;
  wire nn_579, nn_584, nn_561, nwc52, nwc63;
  wire nwc65, nwc66, nwc67, nwc68, nwc69;
  assign overflow = \y[7]_in;
  or eco2 (nn_539, \a[2], \b[2]);
  and eco3 (\y[0], nn_195, nwc66);
  nand eco4 (parity, nn_802, nn_803);
  and eco5 (\y[1], n_508, nwc63);
  and eco6 (\y[2], nn_193, nwc68);
  and eco7 (\y[3], n_492, nwc67);
  and eco8 (\y[4], nn_191, nwc65);
  and eco9 (\y[5], nwc69, nn_190);
  assign \y[6] = \y[7]_in;
  not eco11 (\y[7], nn_69);
  or eco12 (nn_264, wc52, \op[1]);
  or eco13 (nn_475, wc61, \a[5]);
  or eco14 (nn_496, wc42, \a[0]);
  or eco15 (nn_535, \a[4], \b[4]);
  or eco16 (nn_803, nn_451, wc17);
  or eco17 (nn_540, \a[3], \b[3]);
  or eco18 (nn_541, \a[1], \b[1]);
  or eco19 (nn_802, nwc10, nn_195);
  not eco20 (nwc10, nn_451);
  nand eco21 (nn_195, nn_611, nn_612);
  nand eco22 (nn_451, nn_804, nn_805);
  not eco23 (nwc28, nn_551);
  nand eco24 (nn_551, nn_677, nn_678);
  or eco25 (nn_804, nwc12, nn_450);
  not eco26 (nwc12, nn_502);
  nand eco27 (nn_450, nn_811, nn_812);
  nand eco28 (nn_502, nn_806, nn_807);
  or eco29 (nn_805, nn_502, nwc13);
  not eco30 (nwc13, nn_450);
  or eco31 (nn_806, wc20, nn_193);
  or eco32 (nn_193, nwc34, nn_759);
  or eco33 (nn_190, nwc16, nn_729);
  or eco34 (nn_807, nn_190, wc22);
  not eco35 (nwc16, nn_728);
  nand eco36 (nn_729, nn_726, nn_727);
  nand eco37 (nn_728, nn_140, nn_544);
  or eco38 (nn_811, nwc17, nn_191);
  nand eco39 (nn_140, nn_455, nn_475);
  or eco40 (nn_544, nn_696, nwc23);
  not eco41 (nwc17, nn_503);
  or eco42 (nn_191, nwc19, nn_783);
  nand eco43 (nn_503, nn_819, nn_820);
  or eco44 (nn_812, nn_503, wc26);
  or eco45 (nn_726, nwc21, nn_140);
  or eco46 (nn_727, n_725, n_471);
  or eco47 (nn_69, nn_505, nn_264);
  nand eco48 (nn_505, nn_455, nn_705);
  not eco49 (nwc19, nn_782);
  nand eco50 (nn_783, nn_780, n_713);
  nand eco51 (nn_782, n_571, nn_550);
  not eco52 (nwc21, nn_545);
  nand eco53 (nn_545, nn_701, nn_702);
  nand eco54 (nn_696, nn_694, nn_695);
  not eco55 (nwc23, n_472);
  or eco56 (nn_780, nwc28, n_571);
  or eco57 (nn_701, nn_185, nwc31);
  or eco58 (nn_702, nn_264, nn_413);
  or eco59 (nn_550, nn_672, nwc32);
  or eco60 (nn_455, wc7, \b[5]);
  nand eco61 (nn_705, nn_475, nn_413);
  or eco62 (nn_819, wc27, n_508);
  or eco63 (nn_820, n_492, wc21);
  or eco64 (nn_694, nn_185, nn_453);
  or eco65 (nn_695, nn_264, nwc30);
  nand eco66 (nn_413, nn_522, nn_687);
  or eco67 (nn_185, \op[1], \op[0]);
  nand eco68 (nn_453, nn_683, n_710);
  or eco69 (nn_670, nn_264, nwc37);
  not eco70 (nwc30, nn_413);
  not eco71 (nwc31, nn_453);
  nand eco72 (nn_672, nn_670, nn_671);
  not eco73 (nwc32, n_472);
  or eco74 (nn_522, wc3, \b[4]);
  or eco75 (nn_671, nn_185, nn_47);
  nand eco76 (nn_687, n_482, nn_369);
  nand eco77 (nn_683, nn_535, nn_47);
  or eco78 (nn_677, nn_185, nwc38);
  or eco79 (nn_678, nn_264, nn_369);
  nand eco80 (nn_47, nn_662, n_695);
  not eco81 (nwc34, nn_758);
  nand eco82 (nn_759, nn_756, n_668);
  nand eco83 (nn_758, n_565, nn_552);
  not eco84 (nwc37, nn_369);
  nand eco85 (nn_369, n_490, nn_657);
  not eco86 (nwc38, nn_47);
  nand eco87 (nn_410, nn_521, nn_615);
  or eco88 (nn_756, nwc42, n_565);
  or eco89 (nn_552, nn_597, nwc41);
  nand eco90 (nn_657, n_489, nn_410);
  nand eco91 (nn_662, nn_540, nn_56);
  nand eco92 (nn_597, nn_595, nn_596);
  not eco93 (nwc41, n_472);
  not eco94 (nwc42, nn_553);
  nand eco95 (nn_553, nn_602, nn_603);
  nand eco96 (nn_56, nn_620, n_665);
  nand eco97 (nn_611, nn_543, n_471);
  nand eco98 (nn_620, nn_539, nn_41);
  or eco99 (nn_602, nn_185, nwc49);
  or eco100 (nn_603, nn_264, nn_360);
  or eco101 (nn_595, nn_185, nn_41);
  or eco102 (nn_596, nn_264, nwc48);
  or eco103 (nn_521, wc1, \b[2]);
  nand eco104 (nn_615, n_474, nn_360);
  nand eco105 (nn_41, nn_584, n_680);
  or eco106 (nn_612, n_471, n_582);
  not eco107 (nwc48, nn_360);
  nand eco108 (nn_360, n_506, nn_579);
  not eco109 (nwc49, nn_41);
  nand eco110 (nn_543, nn_496, nn_561);
  nand eco111 (nn_579, n_505, nn_496);
  or eco112 (nn_584, nwc52, n_582);
  or eco113 (nn_561, wc47, \b[0]);
  not eco114 (nwc52, nn_541);
  not eco115 (nwc63, nn_69);
  not eco116 (nwc65, nn_69);
  not eco117 (nwc66, nn_69);
  not eco118 (nwc67, nn_69);
  not eco119 (nwc68, nn_69);
  not eco120 (nwc69, nn_69);
endmodule
// cost:141